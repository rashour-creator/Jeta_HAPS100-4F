//##########################################################
// Generated unprefix file for workspace: DW_axi
//##########################################################

`ifdef i_axi___GUARD__DW_AXI_CC_CONSTANTS__VH__
  `define __GUARD__DW_AXI_CC_CONSTANTS__VH__ `i_axi___GUARD__DW_AXI_CC_CONSTANTS__VH__
`endif 

`ifdef i_axi_AXI_USE_RANDOM_SEED
  `define AXI_USE_RANDOM_SEED `i_axi_AXI_USE_RANDOM_SEED
`endif 

`ifdef i_axi_AXI_SEED
  `define AXI_SEED `i_axi_AXI_SEED
`endif 

`ifdef i_axi_USE_FOUNDATION
  `define USE_FOUNDATION `i_axi_USE_FOUNDATION
`endif 

`ifdef i_axi_AXI_DW
  `define AXI_DW `i_axi_AXI_DW
`endif 

`ifdef i_axi_AXI_AW
  `define AXI_AW `i_axi_AXI_AW
`endif 

`ifdef i_axi_AXI_AW_64
  `define AXI_AW_64 `i_axi_AXI_AW_64
`endif 

`ifdef i_axi_AXI_NUM_MASTERS
  `define AXI_NUM_MASTERS `i_axi_AXI_NUM_MASTERS
`endif 

`ifdef i_axi_AXI_NUM_MASTERS_1
  `define AXI_NUM_MASTERS_1 `i_axi_AXI_NUM_MASTERS_1
`endif 

`ifdef i_axi_AXI_HAS_BICMD
  `define AXI_HAS_BICMD `i_axi_AXI_HAS_BICMD
`endif 

`ifdef i_axi_AXI_EN_MULTI_TILE_DLOCK_AVOID
  `define AXI_EN_MULTI_TILE_DLOCK_AVOID `i_axi_AXI_EN_MULTI_TILE_DLOCK_AVOID
`endif 

`ifdef i_axi_AXI_NUM_SYS_MASTERS
  `define AXI_NUM_SYS_MASTERS `i_axi_AXI_NUM_SYS_MASTERS
`endif 

`ifdef i_axi_AXI_NUM_SLAVES
  `define AXI_NUM_SLAVES `i_axi_AXI_NUM_SLAVES
`endif 

`ifdef i_axi_AXI_LOG2_NS
  `define AXI_LOG2_NS `i_axi_AXI_LOG2_NS
`endif 

`ifdef i_axi_AXI_LOG2_NM
  `define AXI_LOG2_NM `i_axi_AXI_LOG2_NM
`endif 

`ifdef i_axi_AXI_LOG2_LCL_NMP1
  `define AXI_LOG2_LCL_NMP1 `i_axi_AXI_LOG2_LCL_NMP1
`endif 

`ifdef i_axi_AXI_LOG2_LCL_NM
  `define AXI_LOG2_LCL_NM `i_axi_AXI_LOG2_LCL_NM
`endif 

`ifdef i_axi_AXI_LOG2_NSP1
  `define AXI_LOG2_NSP1 `i_axi_AXI_LOG2_NSP1
`endif 

`ifdef i_axi_AXI_NSP1
  `define AXI_NSP1 `i_axi_AXI_NSP1
`endif 

`ifdef i_axi_AXI_LOG2_NSP2
  `define AXI_LOG2_NSP2 `i_axi_AXI_LOG2_NSP2
`endif 

`ifdef i_axi_AXI_MIDW
  `define AXI_MIDW `i_axi_AXI_MIDW
`endif 

`ifdef i_axi_AXI_POW2_MIDW
  `define AXI_POW2_MIDW `i_axi_AXI_POW2_MIDW
`endif 

`ifdef i_axi_AXI_SIDW
  `define AXI_SIDW `i_axi_AXI_SIDW
`endif 

`ifdef i_axi_AXI_BLW
  `define AXI_BLW `i_axi_AXI_BLW
`endif 

`ifdef i_axi_AXI_HAS_TZ_SUPPORT
  `define AXI_HAS_TZ_SUPPORT `i_axi_AXI_HAS_TZ_SUPPORT
`endif 

`ifdef i_axi_AXI_TZ_SUPPORT
  `define AXI_TZ_SUPPORT `i_axi_AXI_TZ_SUPPORT
`endif 

`ifdef i_axi_AXI_REMAP_EN
  `define AXI_REMAP_EN `i_axi_AXI_REMAP_EN
`endif 

`ifdef i_axi_AXI_REMAP
  `define AXI_REMAP `i_axi_AXI_REMAP
`endif 

`ifdef i_axi_AXI_HAS_XDCDR
  `define AXI_HAS_XDCDR `i_axi_AXI_HAS_XDCDR
`endif 

`ifdef i_axi_AXI_XDCDR
  `define AXI_XDCDR `i_axi_AXI_XDCDR
`endif 

`ifdef i_axi_AXI_TEST_XDCDR
  `define AXI_TEST_XDCDR `i_axi_AXI_TEST_XDCDR
`endif 

`ifdef i_axi_AXI_INITIAL_LOCKDOWN
  `define AXI_INITIAL_LOCKDOWN `i_axi_AXI_INITIAL_LOCKDOWN
`endif 

`ifdef i_axi_AXI_HAS_LOCKING
  `define AXI_HAS_LOCKING `i_axi_AXI_HAS_LOCKING
`endif 

`ifdef i_axi_AXI_LOCKING
  `define AXI_LOCKING `i_axi_AXI_LOCKING
`endif 

`ifdef i_axi_AXI_LOWPWR_HS_IF
  `define AXI_LOWPWR_HS_IF `i_axi_AXI_LOWPWR_HS_IF
`endif 

`ifdef i_axi_AXI_LOWPWR_NOPX_CNT
  `define AXI_LOWPWR_NOPX_CNT `i_axi_AXI_LOWPWR_NOPX_CNT
`endif 

`ifdef i_axi_AXI_LOG2_LOWPWR_NOPX_CNT
  `define AXI_LOG2_LOWPWR_NOPX_CNT `i_axi_AXI_LOG2_LOWPWR_NOPX_CNT
`endif 

`ifdef i_axi_AXI_INTERFACE_TYPE
  `define AXI_INTERFACE_TYPE `i_axi_AXI_INTERFACE_TYPE
`endif 

`ifdef i_axi_AXI_HAS_AXI4
  `define AXI_HAS_AXI4 `i_axi_AXI_HAS_AXI4
`endif 

`ifdef i_axi_AXI_HAS_QOS
  `define AXI_HAS_QOS `i_axi_AXI_HAS_QOS
`endif 

`ifdef i_axi_AXI_DLOCK_NOTIFY_EN
  `define AXI_DLOCK_NOTIFY_EN `i_axi_AXI_DLOCK_NOTIFY_EN
`endif 

`ifdef i_axi_AXI_DLOCK_TIMEOUT
  `define AXI_DLOCK_TIMEOUT `i_axi_AXI_DLOCK_TIMEOUT
`endif 

`ifdef i_axi_AXI_LOG2_DLOCK_TIMEOUT_P1
  `define AXI_LOG2_DLOCK_TIMEOUT_P1 `i_axi_AXI_LOG2_DLOCK_TIMEOUT_P1
`endif 

`ifdef i_axi_AXI_AR_TMO
  `define AXI_AR_TMO `i_axi_AXI_AR_TMO
`endif 

`ifdef i_axi_AXI_AW_TMO
  `define AXI_AW_TMO `i_axi_AXI_AW_TMO
`endif 

`ifdef i_axi_AXI_W_TMO
  `define AXI_W_TMO `i_axi_AXI_W_TMO
`endif 

`ifdef i_axi_AXI_R_TMO
  `define AXI_R_TMO `i_axi_AXI_R_TMO
`endif 

`ifdef i_axi_AXI_B_TMO
  `define AXI_B_TMO `i_axi_AXI_B_TMO
`endif 

`ifdef i_axi_AXI_AR_PL_ARB
  `define AXI_AR_PL_ARB `i_axi_AXI_AR_PL_ARB
`endif 

`ifdef i_axi_AXI_AW_PL_ARB
  `define AXI_AW_PL_ARB `i_axi_AXI_AW_PL_ARB
`endif 

`ifdef i_axi_AXI_R_PL_ARB
  `define AXI_R_PL_ARB `i_axi_AXI_R_PL_ARB
`endif 

`ifdef i_axi_AXI_W_PL_ARB
  `define AXI_W_PL_ARB `i_axi_AXI_W_PL_ARB
`endif 

`ifdef i_axi_AXI_B_PL_ARB
  `define AXI_B_PL_ARB `i_axi_AXI_B_PL_ARB
`endif 

`ifdef i_axi_AXI_ENCRYPT
  `define AXI_ENCRYPT `i_axi_AXI_ENCRYPT
`endif 

`ifdef i_axi_AXI_MST_PRIORITY_W
  `define AXI_MST_PRIORITY_W `i_axi_AXI_MST_PRIORITY_W
`endif 

`ifdef i_axi_AXI_SLV_PRIORITY_W
  `define AXI_SLV_PRIORITY_W `i_axi_AXI_SLV_PRIORITY_W
`endif 

`ifdef i_axi_AXI_REG_AW_W_PATHS
  `define AXI_REG_AW_W_PATHS `i_axi_AXI_REG_AW_W_PATHS
`endif 

`ifdef i_axi_AXI_MAX_UIDA
  `define AXI_MAX_UIDA `i_axi_AXI_MAX_UIDA
`endif 

`ifdef i_axi_AXI_HAS_LEGAL_ADDR_OVRLP_VAL
  `define AXI_HAS_LEGAL_ADDR_OVRLP_VAL `i_axi_AXI_HAS_LEGAL_ADDR_OVRLP_VAL
`endif 

`ifdef i_axi_AXI_HAS_LEGAL_ADDR_OVRLP
  `define AXI_HAS_LEGAL_ADDR_OVRLP `i_axi_AXI_HAS_LEGAL_ADDR_OVRLP
`endif 

`ifdef i_axi_AXI_VLD_RDY_PARITY_PROT
  `define AXI_VLD_RDY_PARITY_PROT `i_axi_AXI_VLD_RDY_PARITY_PROT
`endif 

`ifdef i_axi_AXI_VLD_RDY_PARITY_MODE
  `define AXI_VLD_RDY_PARITY_MODE `i_axi_AXI_VLD_RDY_PARITY_MODE
`endif 

`ifdef i_axi_AXI_HAS_EVEN_PARITY
  `define AXI_HAS_EVEN_PARITY `i_axi_AXI_HAS_EVEN_PARITY
`endif 

`ifdef i_axi_IFX_RULE_SETUP
  `define IFX_RULE_SETUP `i_axi_IFX_RULE_SETUP
`endif 

`ifdef i_axi_AXI_INTF_PAR_EN
  `define AXI_INTF_PAR_EN `i_axi_AXI_INTF_PAR_EN
`endif 

`ifdef i_axi_AXI_INTF_PARITY_MODE
  `define AXI_INTF_PARITY_MODE `i_axi_AXI_INTF_PARITY_MODE
`endif 

`ifdef i_axi_AXI_MAX_SBW
  `define AXI_MAX_SBW `i_axi_AXI_MAX_SBW
`endif 

`ifdef i_axi_AXI_HAS_AWSB
  `define AXI_HAS_AWSB `i_axi_AXI_HAS_AWSB
`endif 

`ifdef i_axi_AXI_INC_AWSB
  `define AXI_INC_AWSB `i_axi_AXI_INC_AWSB
`endif 

`ifdef i_axi_AXI_AW_SBW
  `define AXI_AW_SBW `i_axi_AXI_AW_SBW
`endif 

`ifdef i_axi_AXI_HAS_WSB
  `define AXI_HAS_WSB `i_axi_AXI_HAS_WSB
`endif 

`ifdef i_axi_AXI_INC_WSB
  `define AXI_INC_WSB `i_axi_AXI_INC_WSB
`endif 

`ifdef i_axi_AXI_W_SBW
  `define AXI_W_SBW `i_axi_AXI_W_SBW
`endif 

`ifdef i_axi_AXI_HAS_BSB
  `define AXI_HAS_BSB `i_axi_AXI_HAS_BSB
`endif 

`ifdef i_axi_AXI_INC_BSB
  `define AXI_INC_BSB `i_axi_AXI_INC_BSB
`endif 

`ifdef i_axi_AXI_B_SBW
  `define AXI_B_SBW `i_axi_AXI_B_SBW
`endif 

`ifdef i_axi_AXI_HAS_ARSB
  `define AXI_HAS_ARSB `i_axi_AXI_HAS_ARSB
`endif 

`ifdef i_axi_AXI_INC_ARSB
  `define AXI_INC_ARSB `i_axi_AXI_INC_ARSB
`endif 

`ifdef i_axi_AXI_AR_SBW
  `define AXI_AR_SBW `i_axi_AXI_AR_SBW
`endif 

`ifdef i_axi_AXI_HAS_RSB
  `define AXI_HAS_RSB `i_axi_AXI_HAS_RSB
`endif 

`ifdef i_axi_AXI_INC_RSB
  `define AXI_INC_RSB `i_axi_AXI_INC_RSB
`endif 

`ifdef i_axi_AXI_R_SBW
  `define AXI_R_SBW `i_axi_AXI_R_SBW
`endif 

`ifdef i_axi_AXI_NV_S0_BY_M1
  `define AXI_NV_S0_BY_M1 `i_axi_AXI_NV_S0_BY_M1
`endif 

`ifdef i_axi_AXI_NV_S0_BY_M2
  `define AXI_NV_S0_BY_M2 `i_axi_AXI_NV_S0_BY_M2
`endif 

`ifdef i_axi_AXI_NV_S0_BY_M3
  `define AXI_NV_S0_BY_M3 `i_axi_AXI_NV_S0_BY_M3
`endif 

`ifdef i_axi_AXI_NV_S0_BY_M4
  `define AXI_NV_S0_BY_M4 `i_axi_AXI_NV_S0_BY_M4
`endif 

`ifdef i_axi_AXI_NV_S0_BY_M5
  `define AXI_NV_S0_BY_M5 `i_axi_AXI_NV_S0_BY_M5
`endif 

`ifdef i_axi_AXI_NV_S0_BY_M6
  `define AXI_NV_S0_BY_M6 `i_axi_AXI_NV_S0_BY_M6
`endif 

`ifdef i_axi_AXI_NV_S0_BY_M7
  `define AXI_NV_S0_BY_M7 `i_axi_AXI_NV_S0_BY_M7
`endif 

`ifdef i_axi_AXI_NV_S0_BY_M8
  `define AXI_NV_S0_BY_M8 `i_axi_AXI_NV_S0_BY_M8
`endif 

`ifdef i_axi_AXI_NV_S0_BY_M9
  `define AXI_NV_S0_BY_M9 `i_axi_AXI_NV_S0_BY_M9
`endif 

`ifdef i_axi_AXI_NV_S0_BY_M10
  `define AXI_NV_S0_BY_M10 `i_axi_AXI_NV_S0_BY_M10
`endif 

`ifdef i_axi_AXI_NV_S0_BY_M11
  `define AXI_NV_S0_BY_M11 `i_axi_AXI_NV_S0_BY_M11
`endif 

`ifdef i_axi_AXI_NV_S0_BY_M12
  `define AXI_NV_S0_BY_M12 `i_axi_AXI_NV_S0_BY_M12
`endif 

`ifdef i_axi_AXI_NV_S0_BY_M13
  `define AXI_NV_S0_BY_M13 `i_axi_AXI_NV_S0_BY_M13
`endif 

`ifdef i_axi_AXI_NV_S0_BY_M14
  `define AXI_NV_S0_BY_M14 `i_axi_AXI_NV_S0_BY_M14
`endif 

`ifdef i_axi_AXI_NV_S0_BY_M15
  `define AXI_NV_S0_BY_M15 `i_axi_AXI_NV_S0_BY_M15
`endif 

`ifdef i_axi_AXI_NV_S0_BY_M16
  `define AXI_NV_S0_BY_M16 `i_axi_AXI_NV_S0_BY_M16
`endif 

`ifdef i_axi_AXI_NV_S1_BY_M1
  `define AXI_NV_S1_BY_M1 `i_axi_AXI_NV_S1_BY_M1
`endif 

`ifdef i_axi_AXI_NV_S1_BY_M2
  `define AXI_NV_S1_BY_M2 `i_axi_AXI_NV_S1_BY_M2
`endif 

`ifdef i_axi_AXI_NV_S1_BY_M3
  `define AXI_NV_S1_BY_M3 `i_axi_AXI_NV_S1_BY_M3
`endif 

`ifdef i_axi_AXI_NV_S1_BY_M4
  `define AXI_NV_S1_BY_M4 `i_axi_AXI_NV_S1_BY_M4
`endif 

`ifdef i_axi_AXI_NV_S1_BY_M5
  `define AXI_NV_S1_BY_M5 `i_axi_AXI_NV_S1_BY_M5
`endif 

`ifdef i_axi_AXI_NV_S1_BY_M6
  `define AXI_NV_S1_BY_M6 `i_axi_AXI_NV_S1_BY_M6
`endif 

`ifdef i_axi_AXI_NV_S1_BY_M7
  `define AXI_NV_S1_BY_M7 `i_axi_AXI_NV_S1_BY_M7
`endif 

`ifdef i_axi_AXI_NV_S1_BY_M8
  `define AXI_NV_S1_BY_M8 `i_axi_AXI_NV_S1_BY_M8
`endif 

`ifdef i_axi_AXI_NV_S1_BY_M9
  `define AXI_NV_S1_BY_M9 `i_axi_AXI_NV_S1_BY_M9
`endif 

`ifdef i_axi_AXI_NV_S1_BY_M10
  `define AXI_NV_S1_BY_M10 `i_axi_AXI_NV_S1_BY_M10
`endif 

`ifdef i_axi_AXI_NV_S1_BY_M11
  `define AXI_NV_S1_BY_M11 `i_axi_AXI_NV_S1_BY_M11
`endif 

`ifdef i_axi_AXI_NV_S1_BY_M12
  `define AXI_NV_S1_BY_M12 `i_axi_AXI_NV_S1_BY_M12
`endif 

`ifdef i_axi_AXI_NV_S1_BY_M13
  `define AXI_NV_S1_BY_M13 `i_axi_AXI_NV_S1_BY_M13
`endif 

`ifdef i_axi_AXI_NV_S1_BY_M14
  `define AXI_NV_S1_BY_M14 `i_axi_AXI_NV_S1_BY_M14
`endif 

`ifdef i_axi_AXI_NV_S1_BY_M15
  `define AXI_NV_S1_BY_M15 `i_axi_AXI_NV_S1_BY_M15
`endif 

`ifdef i_axi_AXI_NV_S1_BY_M16
  `define AXI_NV_S1_BY_M16 `i_axi_AXI_NV_S1_BY_M16
`endif 

`ifdef i_axi_AXI_NV_S2_BY_M1
  `define AXI_NV_S2_BY_M1 `i_axi_AXI_NV_S2_BY_M1
`endif 

`ifdef i_axi_AXI_NV_S2_BY_M2
  `define AXI_NV_S2_BY_M2 `i_axi_AXI_NV_S2_BY_M2
`endif 

`ifdef i_axi_AXI_NV_S2_BY_M3
  `define AXI_NV_S2_BY_M3 `i_axi_AXI_NV_S2_BY_M3
`endif 

`ifdef i_axi_AXI_NV_S2_BY_M4
  `define AXI_NV_S2_BY_M4 `i_axi_AXI_NV_S2_BY_M4
`endif 

`ifdef i_axi_AXI_NV_S2_BY_M5
  `define AXI_NV_S2_BY_M5 `i_axi_AXI_NV_S2_BY_M5
`endif 

`ifdef i_axi_AXI_NV_S2_BY_M6
  `define AXI_NV_S2_BY_M6 `i_axi_AXI_NV_S2_BY_M6
`endif 

`ifdef i_axi_AXI_NV_S2_BY_M7
  `define AXI_NV_S2_BY_M7 `i_axi_AXI_NV_S2_BY_M7
`endif 

`ifdef i_axi_AXI_NV_S2_BY_M8
  `define AXI_NV_S2_BY_M8 `i_axi_AXI_NV_S2_BY_M8
`endif 

`ifdef i_axi_AXI_NV_S2_BY_M9
  `define AXI_NV_S2_BY_M9 `i_axi_AXI_NV_S2_BY_M9
`endif 

`ifdef i_axi_AXI_NV_S2_BY_M10
  `define AXI_NV_S2_BY_M10 `i_axi_AXI_NV_S2_BY_M10
`endif 

`ifdef i_axi_AXI_NV_S2_BY_M11
  `define AXI_NV_S2_BY_M11 `i_axi_AXI_NV_S2_BY_M11
`endif 

`ifdef i_axi_AXI_NV_S2_BY_M12
  `define AXI_NV_S2_BY_M12 `i_axi_AXI_NV_S2_BY_M12
`endif 

`ifdef i_axi_AXI_NV_S2_BY_M13
  `define AXI_NV_S2_BY_M13 `i_axi_AXI_NV_S2_BY_M13
`endif 

`ifdef i_axi_AXI_NV_S2_BY_M14
  `define AXI_NV_S2_BY_M14 `i_axi_AXI_NV_S2_BY_M14
`endif 

`ifdef i_axi_AXI_NV_S2_BY_M15
  `define AXI_NV_S2_BY_M15 `i_axi_AXI_NV_S2_BY_M15
`endif 

`ifdef i_axi_AXI_NV_S2_BY_M16
  `define AXI_NV_S2_BY_M16 `i_axi_AXI_NV_S2_BY_M16
`endif 

`ifdef i_axi_AXI_NV_S3_BY_M1
  `define AXI_NV_S3_BY_M1 `i_axi_AXI_NV_S3_BY_M1
`endif 

`ifdef i_axi_AXI_NV_S3_BY_M2
  `define AXI_NV_S3_BY_M2 `i_axi_AXI_NV_S3_BY_M2
`endif 

`ifdef i_axi_AXI_NV_S3_BY_M3
  `define AXI_NV_S3_BY_M3 `i_axi_AXI_NV_S3_BY_M3
`endif 

`ifdef i_axi_AXI_NV_S3_BY_M4
  `define AXI_NV_S3_BY_M4 `i_axi_AXI_NV_S3_BY_M4
`endif 

`ifdef i_axi_AXI_NV_S3_BY_M5
  `define AXI_NV_S3_BY_M5 `i_axi_AXI_NV_S3_BY_M5
`endif 

`ifdef i_axi_AXI_NV_S3_BY_M6
  `define AXI_NV_S3_BY_M6 `i_axi_AXI_NV_S3_BY_M6
`endif 

`ifdef i_axi_AXI_NV_S3_BY_M7
  `define AXI_NV_S3_BY_M7 `i_axi_AXI_NV_S3_BY_M7
`endif 

`ifdef i_axi_AXI_NV_S3_BY_M8
  `define AXI_NV_S3_BY_M8 `i_axi_AXI_NV_S3_BY_M8
`endif 

`ifdef i_axi_AXI_NV_S3_BY_M9
  `define AXI_NV_S3_BY_M9 `i_axi_AXI_NV_S3_BY_M9
`endif 

`ifdef i_axi_AXI_NV_S3_BY_M10
  `define AXI_NV_S3_BY_M10 `i_axi_AXI_NV_S3_BY_M10
`endif 

`ifdef i_axi_AXI_NV_S3_BY_M11
  `define AXI_NV_S3_BY_M11 `i_axi_AXI_NV_S3_BY_M11
`endif 

`ifdef i_axi_AXI_NV_S3_BY_M12
  `define AXI_NV_S3_BY_M12 `i_axi_AXI_NV_S3_BY_M12
`endif 

`ifdef i_axi_AXI_NV_S3_BY_M13
  `define AXI_NV_S3_BY_M13 `i_axi_AXI_NV_S3_BY_M13
`endif 

`ifdef i_axi_AXI_NV_S3_BY_M14
  `define AXI_NV_S3_BY_M14 `i_axi_AXI_NV_S3_BY_M14
`endif 

`ifdef i_axi_AXI_NV_S3_BY_M15
  `define AXI_NV_S3_BY_M15 `i_axi_AXI_NV_S3_BY_M15
`endif 

`ifdef i_axi_AXI_NV_S3_BY_M16
  `define AXI_NV_S3_BY_M16 `i_axi_AXI_NV_S3_BY_M16
`endif 

`ifdef i_axi_AXI_NV_S4_BY_M1
  `define AXI_NV_S4_BY_M1 `i_axi_AXI_NV_S4_BY_M1
`endif 

`ifdef i_axi_AXI_NV_S4_BY_M2
  `define AXI_NV_S4_BY_M2 `i_axi_AXI_NV_S4_BY_M2
`endif 

`ifdef i_axi_AXI_NV_S4_BY_M3
  `define AXI_NV_S4_BY_M3 `i_axi_AXI_NV_S4_BY_M3
`endif 

`ifdef i_axi_AXI_NV_S4_BY_M4
  `define AXI_NV_S4_BY_M4 `i_axi_AXI_NV_S4_BY_M4
`endif 

`ifdef i_axi_AXI_NV_S4_BY_M5
  `define AXI_NV_S4_BY_M5 `i_axi_AXI_NV_S4_BY_M5
`endif 

`ifdef i_axi_AXI_NV_S4_BY_M6
  `define AXI_NV_S4_BY_M6 `i_axi_AXI_NV_S4_BY_M6
`endif 

`ifdef i_axi_AXI_NV_S4_BY_M7
  `define AXI_NV_S4_BY_M7 `i_axi_AXI_NV_S4_BY_M7
`endif 

`ifdef i_axi_AXI_NV_S4_BY_M8
  `define AXI_NV_S4_BY_M8 `i_axi_AXI_NV_S4_BY_M8
`endif 

`ifdef i_axi_AXI_NV_S4_BY_M9
  `define AXI_NV_S4_BY_M9 `i_axi_AXI_NV_S4_BY_M9
`endif 

`ifdef i_axi_AXI_NV_S4_BY_M10
  `define AXI_NV_S4_BY_M10 `i_axi_AXI_NV_S4_BY_M10
`endif 

`ifdef i_axi_AXI_NV_S4_BY_M11
  `define AXI_NV_S4_BY_M11 `i_axi_AXI_NV_S4_BY_M11
`endif 

`ifdef i_axi_AXI_NV_S4_BY_M12
  `define AXI_NV_S4_BY_M12 `i_axi_AXI_NV_S4_BY_M12
`endif 

`ifdef i_axi_AXI_NV_S4_BY_M13
  `define AXI_NV_S4_BY_M13 `i_axi_AXI_NV_S4_BY_M13
`endif 

`ifdef i_axi_AXI_NV_S4_BY_M14
  `define AXI_NV_S4_BY_M14 `i_axi_AXI_NV_S4_BY_M14
`endif 

`ifdef i_axi_AXI_NV_S4_BY_M15
  `define AXI_NV_S4_BY_M15 `i_axi_AXI_NV_S4_BY_M15
`endif 

`ifdef i_axi_AXI_NV_S4_BY_M16
  `define AXI_NV_S4_BY_M16 `i_axi_AXI_NV_S4_BY_M16
`endif 

`ifdef i_axi_AXI_NV_S5_BY_M1
  `define AXI_NV_S5_BY_M1 `i_axi_AXI_NV_S5_BY_M1
`endif 

`ifdef i_axi_AXI_NV_S5_BY_M2
  `define AXI_NV_S5_BY_M2 `i_axi_AXI_NV_S5_BY_M2
`endif 

`ifdef i_axi_AXI_NV_S5_BY_M3
  `define AXI_NV_S5_BY_M3 `i_axi_AXI_NV_S5_BY_M3
`endif 

`ifdef i_axi_AXI_NV_S5_BY_M4
  `define AXI_NV_S5_BY_M4 `i_axi_AXI_NV_S5_BY_M4
`endif 

`ifdef i_axi_AXI_NV_S5_BY_M5
  `define AXI_NV_S5_BY_M5 `i_axi_AXI_NV_S5_BY_M5
`endif 

`ifdef i_axi_AXI_NV_S5_BY_M6
  `define AXI_NV_S5_BY_M6 `i_axi_AXI_NV_S5_BY_M6
`endif 

`ifdef i_axi_AXI_NV_S5_BY_M7
  `define AXI_NV_S5_BY_M7 `i_axi_AXI_NV_S5_BY_M7
`endif 

`ifdef i_axi_AXI_NV_S5_BY_M8
  `define AXI_NV_S5_BY_M8 `i_axi_AXI_NV_S5_BY_M8
`endif 

`ifdef i_axi_AXI_NV_S5_BY_M9
  `define AXI_NV_S5_BY_M9 `i_axi_AXI_NV_S5_BY_M9
`endif 

`ifdef i_axi_AXI_NV_S5_BY_M10
  `define AXI_NV_S5_BY_M10 `i_axi_AXI_NV_S5_BY_M10
`endif 

`ifdef i_axi_AXI_NV_S5_BY_M11
  `define AXI_NV_S5_BY_M11 `i_axi_AXI_NV_S5_BY_M11
`endif 

`ifdef i_axi_AXI_NV_S5_BY_M12
  `define AXI_NV_S5_BY_M12 `i_axi_AXI_NV_S5_BY_M12
`endif 

`ifdef i_axi_AXI_NV_S5_BY_M13
  `define AXI_NV_S5_BY_M13 `i_axi_AXI_NV_S5_BY_M13
`endif 

`ifdef i_axi_AXI_NV_S5_BY_M14
  `define AXI_NV_S5_BY_M14 `i_axi_AXI_NV_S5_BY_M14
`endif 

`ifdef i_axi_AXI_NV_S5_BY_M15
  `define AXI_NV_S5_BY_M15 `i_axi_AXI_NV_S5_BY_M15
`endif 

`ifdef i_axi_AXI_NV_S5_BY_M16
  `define AXI_NV_S5_BY_M16 `i_axi_AXI_NV_S5_BY_M16
`endif 

`ifdef i_axi_AXI_NV_S6_BY_M1
  `define AXI_NV_S6_BY_M1 `i_axi_AXI_NV_S6_BY_M1
`endif 

`ifdef i_axi_AXI_NV_S6_BY_M2
  `define AXI_NV_S6_BY_M2 `i_axi_AXI_NV_S6_BY_M2
`endif 

`ifdef i_axi_AXI_NV_S6_BY_M3
  `define AXI_NV_S6_BY_M3 `i_axi_AXI_NV_S6_BY_M3
`endif 

`ifdef i_axi_AXI_NV_S6_BY_M4
  `define AXI_NV_S6_BY_M4 `i_axi_AXI_NV_S6_BY_M4
`endif 

`ifdef i_axi_AXI_NV_S6_BY_M5
  `define AXI_NV_S6_BY_M5 `i_axi_AXI_NV_S6_BY_M5
`endif 

`ifdef i_axi_AXI_NV_S6_BY_M6
  `define AXI_NV_S6_BY_M6 `i_axi_AXI_NV_S6_BY_M6
`endif 

`ifdef i_axi_AXI_NV_S6_BY_M7
  `define AXI_NV_S6_BY_M7 `i_axi_AXI_NV_S6_BY_M7
`endif 

`ifdef i_axi_AXI_NV_S6_BY_M8
  `define AXI_NV_S6_BY_M8 `i_axi_AXI_NV_S6_BY_M8
`endif 

`ifdef i_axi_AXI_NV_S6_BY_M9
  `define AXI_NV_S6_BY_M9 `i_axi_AXI_NV_S6_BY_M9
`endif 

`ifdef i_axi_AXI_NV_S6_BY_M10
  `define AXI_NV_S6_BY_M10 `i_axi_AXI_NV_S6_BY_M10
`endif 

`ifdef i_axi_AXI_NV_S6_BY_M11
  `define AXI_NV_S6_BY_M11 `i_axi_AXI_NV_S6_BY_M11
`endif 

`ifdef i_axi_AXI_NV_S6_BY_M12
  `define AXI_NV_S6_BY_M12 `i_axi_AXI_NV_S6_BY_M12
`endif 

`ifdef i_axi_AXI_NV_S6_BY_M13
  `define AXI_NV_S6_BY_M13 `i_axi_AXI_NV_S6_BY_M13
`endif 

`ifdef i_axi_AXI_NV_S6_BY_M14
  `define AXI_NV_S6_BY_M14 `i_axi_AXI_NV_S6_BY_M14
`endif 

`ifdef i_axi_AXI_NV_S6_BY_M15
  `define AXI_NV_S6_BY_M15 `i_axi_AXI_NV_S6_BY_M15
`endif 

`ifdef i_axi_AXI_NV_S6_BY_M16
  `define AXI_NV_S6_BY_M16 `i_axi_AXI_NV_S6_BY_M16
`endif 

`ifdef i_axi_AXI_NV_S7_BY_M1
  `define AXI_NV_S7_BY_M1 `i_axi_AXI_NV_S7_BY_M1
`endif 

`ifdef i_axi_AXI_NV_S7_BY_M2
  `define AXI_NV_S7_BY_M2 `i_axi_AXI_NV_S7_BY_M2
`endif 

`ifdef i_axi_AXI_NV_S7_BY_M3
  `define AXI_NV_S7_BY_M3 `i_axi_AXI_NV_S7_BY_M3
`endif 

`ifdef i_axi_AXI_NV_S7_BY_M4
  `define AXI_NV_S7_BY_M4 `i_axi_AXI_NV_S7_BY_M4
`endif 

`ifdef i_axi_AXI_NV_S7_BY_M5
  `define AXI_NV_S7_BY_M5 `i_axi_AXI_NV_S7_BY_M5
`endif 

`ifdef i_axi_AXI_NV_S7_BY_M6
  `define AXI_NV_S7_BY_M6 `i_axi_AXI_NV_S7_BY_M6
`endif 

`ifdef i_axi_AXI_NV_S7_BY_M7
  `define AXI_NV_S7_BY_M7 `i_axi_AXI_NV_S7_BY_M7
`endif 

`ifdef i_axi_AXI_NV_S7_BY_M8
  `define AXI_NV_S7_BY_M8 `i_axi_AXI_NV_S7_BY_M8
`endif 

`ifdef i_axi_AXI_NV_S7_BY_M9
  `define AXI_NV_S7_BY_M9 `i_axi_AXI_NV_S7_BY_M9
`endif 

`ifdef i_axi_AXI_NV_S7_BY_M10
  `define AXI_NV_S7_BY_M10 `i_axi_AXI_NV_S7_BY_M10
`endif 

`ifdef i_axi_AXI_NV_S7_BY_M11
  `define AXI_NV_S7_BY_M11 `i_axi_AXI_NV_S7_BY_M11
`endif 

`ifdef i_axi_AXI_NV_S7_BY_M12
  `define AXI_NV_S7_BY_M12 `i_axi_AXI_NV_S7_BY_M12
`endif 

`ifdef i_axi_AXI_NV_S7_BY_M13
  `define AXI_NV_S7_BY_M13 `i_axi_AXI_NV_S7_BY_M13
`endif 

`ifdef i_axi_AXI_NV_S7_BY_M14
  `define AXI_NV_S7_BY_M14 `i_axi_AXI_NV_S7_BY_M14
`endif 

`ifdef i_axi_AXI_NV_S7_BY_M15
  `define AXI_NV_S7_BY_M15 `i_axi_AXI_NV_S7_BY_M15
`endif 

`ifdef i_axi_AXI_NV_S7_BY_M16
  `define AXI_NV_S7_BY_M16 `i_axi_AXI_NV_S7_BY_M16
`endif 

`ifdef i_axi_AXI_NV_S8_BY_M1
  `define AXI_NV_S8_BY_M1 `i_axi_AXI_NV_S8_BY_M1
`endif 

`ifdef i_axi_AXI_NV_S8_BY_M2
  `define AXI_NV_S8_BY_M2 `i_axi_AXI_NV_S8_BY_M2
`endif 

`ifdef i_axi_AXI_NV_S8_BY_M3
  `define AXI_NV_S8_BY_M3 `i_axi_AXI_NV_S8_BY_M3
`endif 

`ifdef i_axi_AXI_NV_S8_BY_M4
  `define AXI_NV_S8_BY_M4 `i_axi_AXI_NV_S8_BY_M4
`endif 

`ifdef i_axi_AXI_NV_S8_BY_M5
  `define AXI_NV_S8_BY_M5 `i_axi_AXI_NV_S8_BY_M5
`endif 

`ifdef i_axi_AXI_NV_S8_BY_M6
  `define AXI_NV_S8_BY_M6 `i_axi_AXI_NV_S8_BY_M6
`endif 

`ifdef i_axi_AXI_NV_S8_BY_M7
  `define AXI_NV_S8_BY_M7 `i_axi_AXI_NV_S8_BY_M7
`endif 

`ifdef i_axi_AXI_NV_S8_BY_M8
  `define AXI_NV_S8_BY_M8 `i_axi_AXI_NV_S8_BY_M8
`endif 

`ifdef i_axi_AXI_NV_S8_BY_M9
  `define AXI_NV_S8_BY_M9 `i_axi_AXI_NV_S8_BY_M9
`endif 

`ifdef i_axi_AXI_NV_S8_BY_M10
  `define AXI_NV_S8_BY_M10 `i_axi_AXI_NV_S8_BY_M10
`endif 

`ifdef i_axi_AXI_NV_S8_BY_M11
  `define AXI_NV_S8_BY_M11 `i_axi_AXI_NV_S8_BY_M11
`endif 

`ifdef i_axi_AXI_NV_S8_BY_M12
  `define AXI_NV_S8_BY_M12 `i_axi_AXI_NV_S8_BY_M12
`endif 

`ifdef i_axi_AXI_NV_S8_BY_M13
  `define AXI_NV_S8_BY_M13 `i_axi_AXI_NV_S8_BY_M13
`endif 

`ifdef i_axi_AXI_NV_S8_BY_M14
  `define AXI_NV_S8_BY_M14 `i_axi_AXI_NV_S8_BY_M14
`endif 

`ifdef i_axi_AXI_NV_S8_BY_M15
  `define AXI_NV_S8_BY_M15 `i_axi_AXI_NV_S8_BY_M15
`endif 

`ifdef i_axi_AXI_NV_S8_BY_M16
  `define AXI_NV_S8_BY_M16 `i_axi_AXI_NV_S8_BY_M16
`endif 

`ifdef i_axi_AXI_NV_S9_BY_M1
  `define AXI_NV_S9_BY_M1 `i_axi_AXI_NV_S9_BY_M1
`endif 

`ifdef i_axi_AXI_NV_S9_BY_M2
  `define AXI_NV_S9_BY_M2 `i_axi_AXI_NV_S9_BY_M2
`endif 

`ifdef i_axi_AXI_NV_S9_BY_M3
  `define AXI_NV_S9_BY_M3 `i_axi_AXI_NV_S9_BY_M3
`endif 

`ifdef i_axi_AXI_NV_S9_BY_M4
  `define AXI_NV_S9_BY_M4 `i_axi_AXI_NV_S9_BY_M4
`endif 

`ifdef i_axi_AXI_NV_S9_BY_M5
  `define AXI_NV_S9_BY_M5 `i_axi_AXI_NV_S9_BY_M5
`endif 

`ifdef i_axi_AXI_NV_S9_BY_M6
  `define AXI_NV_S9_BY_M6 `i_axi_AXI_NV_S9_BY_M6
`endif 

`ifdef i_axi_AXI_NV_S9_BY_M7
  `define AXI_NV_S9_BY_M7 `i_axi_AXI_NV_S9_BY_M7
`endif 

`ifdef i_axi_AXI_NV_S9_BY_M8
  `define AXI_NV_S9_BY_M8 `i_axi_AXI_NV_S9_BY_M8
`endif 

`ifdef i_axi_AXI_NV_S9_BY_M9
  `define AXI_NV_S9_BY_M9 `i_axi_AXI_NV_S9_BY_M9
`endif 

`ifdef i_axi_AXI_NV_S9_BY_M10
  `define AXI_NV_S9_BY_M10 `i_axi_AXI_NV_S9_BY_M10
`endif 

`ifdef i_axi_AXI_NV_S9_BY_M11
  `define AXI_NV_S9_BY_M11 `i_axi_AXI_NV_S9_BY_M11
`endif 

`ifdef i_axi_AXI_NV_S9_BY_M12
  `define AXI_NV_S9_BY_M12 `i_axi_AXI_NV_S9_BY_M12
`endif 

`ifdef i_axi_AXI_NV_S9_BY_M13
  `define AXI_NV_S9_BY_M13 `i_axi_AXI_NV_S9_BY_M13
`endif 

`ifdef i_axi_AXI_NV_S9_BY_M14
  `define AXI_NV_S9_BY_M14 `i_axi_AXI_NV_S9_BY_M14
`endif 

`ifdef i_axi_AXI_NV_S9_BY_M15
  `define AXI_NV_S9_BY_M15 `i_axi_AXI_NV_S9_BY_M15
`endif 

`ifdef i_axi_AXI_NV_S9_BY_M16
  `define AXI_NV_S9_BY_M16 `i_axi_AXI_NV_S9_BY_M16
`endif 

`ifdef i_axi_AXI_NV_S10_BY_M1
  `define AXI_NV_S10_BY_M1 `i_axi_AXI_NV_S10_BY_M1
`endif 

`ifdef i_axi_AXI_NV_S10_BY_M2
  `define AXI_NV_S10_BY_M2 `i_axi_AXI_NV_S10_BY_M2
`endif 

`ifdef i_axi_AXI_NV_S10_BY_M3
  `define AXI_NV_S10_BY_M3 `i_axi_AXI_NV_S10_BY_M3
`endif 

`ifdef i_axi_AXI_NV_S10_BY_M4
  `define AXI_NV_S10_BY_M4 `i_axi_AXI_NV_S10_BY_M4
`endif 

`ifdef i_axi_AXI_NV_S10_BY_M5
  `define AXI_NV_S10_BY_M5 `i_axi_AXI_NV_S10_BY_M5
`endif 

`ifdef i_axi_AXI_NV_S10_BY_M6
  `define AXI_NV_S10_BY_M6 `i_axi_AXI_NV_S10_BY_M6
`endif 

`ifdef i_axi_AXI_NV_S10_BY_M7
  `define AXI_NV_S10_BY_M7 `i_axi_AXI_NV_S10_BY_M7
`endif 

`ifdef i_axi_AXI_NV_S10_BY_M8
  `define AXI_NV_S10_BY_M8 `i_axi_AXI_NV_S10_BY_M8
`endif 

`ifdef i_axi_AXI_NV_S10_BY_M9
  `define AXI_NV_S10_BY_M9 `i_axi_AXI_NV_S10_BY_M9
`endif 

`ifdef i_axi_AXI_NV_S10_BY_M10
  `define AXI_NV_S10_BY_M10 `i_axi_AXI_NV_S10_BY_M10
`endif 

`ifdef i_axi_AXI_NV_S10_BY_M11
  `define AXI_NV_S10_BY_M11 `i_axi_AXI_NV_S10_BY_M11
`endif 

`ifdef i_axi_AXI_NV_S10_BY_M12
  `define AXI_NV_S10_BY_M12 `i_axi_AXI_NV_S10_BY_M12
`endif 

`ifdef i_axi_AXI_NV_S10_BY_M13
  `define AXI_NV_S10_BY_M13 `i_axi_AXI_NV_S10_BY_M13
`endif 

`ifdef i_axi_AXI_NV_S10_BY_M14
  `define AXI_NV_S10_BY_M14 `i_axi_AXI_NV_S10_BY_M14
`endif 

`ifdef i_axi_AXI_NV_S10_BY_M15
  `define AXI_NV_S10_BY_M15 `i_axi_AXI_NV_S10_BY_M15
`endif 

`ifdef i_axi_AXI_NV_S10_BY_M16
  `define AXI_NV_S10_BY_M16 `i_axi_AXI_NV_S10_BY_M16
`endif 

`ifdef i_axi_AXI_NV_S11_BY_M1
  `define AXI_NV_S11_BY_M1 `i_axi_AXI_NV_S11_BY_M1
`endif 

`ifdef i_axi_AXI_NV_S11_BY_M2
  `define AXI_NV_S11_BY_M2 `i_axi_AXI_NV_S11_BY_M2
`endif 

`ifdef i_axi_AXI_NV_S11_BY_M3
  `define AXI_NV_S11_BY_M3 `i_axi_AXI_NV_S11_BY_M3
`endif 

`ifdef i_axi_AXI_NV_S11_BY_M4
  `define AXI_NV_S11_BY_M4 `i_axi_AXI_NV_S11_BY_M4
`endif 

`ifdef i_axi_AXI_NV_S11_BY_M5
  `define AXI_NV_S11_BY_M5 `i_axi_AXI_NV_S11_BY_M5
`endif 

`ifdef i_axi_AXI_NV_S11_BY_M6
  `define AXI_NV_S11_BY_M6 `i_axi_AXI_NV_S11_BY_M6
`endif 

`ifdef i_axi_AXI_NV_S11_BY_M7
  `define AXI_NV_S11_BY_M7 `i_axi_AXI_NV_S11_BY_M7
`endif 

`ifdef i_axi_AXI_NV_S11_BY_M8
  `define AXI_NV_S11_BY_M8 `i_axi_AXI_NV_S11_BY_M8
`endif 

`ifdef i_axi_AXI_NV_S11_BY_M9
  `define AXI_NV_S11_BY_M9 `i_axi_AXI_NV_S11_BY_M9
`endif 

`ifdef i_axi_AXI_NV_S11_BY_M10
  `define AXI_NV_S11_BY_M10 `i_axi_AXI_NV_S11_BY_M10
`endif 

`ifdef i_axi_AXI_NV_S11_BY_M11
  `define AXI_NV_S11_BY_M11 `i_axi_AXI_NV_S11_BY_M11
`endif 

`ifdef i_axi_AXI_NV_S11_BY_M12
  `define AXI_NV_S11_BY_M12 `i_axi_AXI_NV_S11_BY_M12
`endif 

`ifdef i_axi_AXI_NV_S11_BY_M13
  `define AXI_NV_S11_BY_M13 `i_axi_AXI_NV_S11_BY_M13
`endif 

`ifdef i_axi_AXI_NV_S11_BY_M14
  `define AXI_NV_S11_BY_M14 `i_axi_AXI_NV_S11_BY_M14
`endif 

`ifdef i_axi_AXI_NV_S11_BY_M15
  `define AXI_NV_S11_BY_M15 `i_axi_AXI_NV_S11_BY_M15
`endif 

`ifdef i_axi_AXI_NV_S11_BY_M16
  `define AXI_NV_S11_BY_M16 `i_axi_AXI_NV_S11_BY_M16
`endif 

`ifdef i_axi_AXI_NV_S12_BY_M1
  `define AXI_NV_S12_BY_M1 `i_axi_AXI_NV_S12_BY_M1
`endif 

`ifdef i_axi_AXI_NV_S12_BY_M2
  `define AXI_NV_S12_BY_M2 `i_axi_AXI_NV_S12_BY_M2
`endif 

`ifdef i_axi_AXI_NV_S12_BY_M3
  `define AXI_NV_S12_BY_M3 `i_axi_AXI_NV_S12_BY_M3
`endif 

`ifdef i_axi_AXI_NV_S12_BY_M4
  `define AXI_NV_S12_BY_M4 `i_axi_AXI_NV_S12_BY_M4
`endif 

`ifdef i_axi_AXI_NV_S12_BY_M5
  `define AXI_NV_S12_BY_M5 `i_axi_AXI_NV_S12_BY_M5
`endif 

`ifdef i_axi_AXI_NV_S12_BY_M6
  `define AXI_NV_S12_BY_M6 `i_axi_AXI_NV_S12_BY_M6
`endif 

`ifdef i_axi_AXI_NV_S12_BY_M7
  `define AXI_NV_S12_BY_M7 `i_axi_AXI_NV_S12_BY_M7
`endif 

`ifdef i_axi_AXI_NV_S12_BY_M8
  `define AXI_NV_S12_BY_M8 `i_axi_AXI_NV_S12_BY_M8
`endif 

`ifdef i_axi_AXI_NV_S12_BY_M9
  `define AXI_NV_S12_BY_M9 `i_axi_AXI_NV_S12_BY_M9
`endif 

`ifdef i_axi_AXI_NV_S12_BY_M10
  `define AXI_NV_S12_BY_M10 `i_axi_AXI_NV_S12_BY_M10
`endif 

`ifdef i_axi_AXI_NV_S12_BY_M11
  `define AXI_NV_S12_BY_M11 `i_axi_AXI_NV_S12_BY_M11
`endif 

`ifdef i_axi_AXI_NV_S12_BY_M12
  `define AXI_NV_S12_BY_M12 `i_axi_AXI_NV_S12_BY_M12
`endif 

`ifdef i_axi_AXI_NV_S12_BY_M13
  `define AXI_NV_S12_BY_M13 `i_axi_AXI_NV_S12_BY_M13
`endif 

`ifdef i_axi_AXI_NV_S12_BY_M14
  `define AXI_NV_S12_BY_M14 `i_axi_AXI_NV_S12_BY_M14
`endif 

`ifdef i_axi_AXI_NV_S12_BY_M15
  `define AXI_NV_S12_BY_M15 `i_axi_AXI_NV_S12_BY_M15
`endif 

`ifdef i_axi_AXI_NV_S12_BY_M16
  `define AXI_NV_S12_BY_M16 `i_axi_AXI_NV_S12_BY_M16
`endif 

`ifdef i_axi_AXI_NV_S13_BY_M1
  `define AXI_NV_S13_BY_M1 `i_axi_AXI_NV_S13_BY_M1
`endif 

`ifdef i_axi_AXI_NV_S13_BY_M2
  `define AXI_NV_S13_BY_M2 `i_axi_AXI_NV_S13_BY_M2
`endif 

`ifdef i_axi_AXI_NV_S13_BY_M3
  `define AXI_NV_S13_BY_M3 `i_axi_AXI_NV_S13_BY_M3
`endif 

`ifdef i_axi_AXI_NV_S13_BY_M4
  `define AXI_NV_S13_BY_M4 `i_axi_AXI_NV_S13_BY_M4
`endif 

`ifdef i_axi_AXI_NV_S13_BY_M5
  `define AXI_NV_S13_BY_M5 `i_axi_AXI_NV_S13_BY_M5
`endif 

`ifdef i_axi_AXI_NV_S13_BY_M6
  `define AXI_NV_S13_BY_M6 `i_axi_AXI_NV_S13_BY_M6
`endif 

`ifdef i_axi_AXI_NV_S13_BY_M7
  `define AXI_NV_S13_BY_M7 `i_axi_AXI_NV_S13_BY_M7
`endif 

`ifdef i_axi_AXI_NV_S13_BY_M8
  `define AXI_NV_S13_BY_M8 `i_axi_AXI_NV_S13_BY_M8
`endif 

`ifdef i_axi_AXI_NV_S13_BY_M9
  `define AXI_NV_S13_BY_M9 `i_axi_AXI_NV_S13_BY_M9
`endif 

`ifdef i_axi_AXI_NV_S13_BY_M10
  `define AXI_NV_S13_BY_M10 `i_axi_AXI_NV_S13_BY_M10
`endif 

`ifdef i_axi_AXI_NV_S13_BY_M11
  `define AXI_NV_S13_BY_M11 `i_axi_AXI_NV_S13_BY_M11
`endif 

`ifdef i_axi_AXI_NV_S13_BY_M12
  `define AXI_NV_S13_BY_M12 `i_axi_AXI_NV_S13_BY_M12
`endif 

`ifdef i_axi_AXI_NV_S13_BY_M13
  `define AXI_NV_S13_BY_M13 `i_axi_AXI_NV_S13_BY_M13
`endif 

`ifdef i_axi_AXI_NV_S13_BY_M14
  `define AXI_NV_S13_BY_M14 `i_axi_AXI_NV_S13_BY_M14
`endif 

`ifdef i_axi_AXI_NV_S13_BY_M15
  `define AXI_NV_S13_BY_M15 `i_axi_AXI_NV_S13_BY_M15
`endif 

`ifdef i_axi_AXI_NV_S13_BY_M16
  `define AXI_NV_S13_BY_M16 `i_axi_AXI_NV_S13_BY_M16
`endif 

`ifdef i_axi_AXI_NV_S14_BY_M1
  `define AXI_NV_S14_BY_M1 `i_axi_AXI_NV_S14_BY_M1
`endif 

`ifdef i_axi_AXI_NV_S14_BY_M2
  `define AXI_NV_S14_BY_M2 `i_axi_AXI_NV_S14_BY_M2
`endif 

`ifdef i_axi_AXI_NV_S14_BY_M3
  `define AXI_NV_S14_BY_M3 `i_axi_AXI_NV_S14_BY_M3
`endif 

`ifdef i_axi_AXI_NV_S14_BY_M4
  `define AXI_NV_S14_BY_M4 `i_axi_AXI_NV_S14_BY_M4
`endif 

`ifdef i_axi_AXI_NV_S14_BY_M5
  `define AXI_NV_S14_BY_M5 `i_axi_AXI_NV_S14_BY_M5
`endif 

`ifdef i_axi_AXI_NV_S14_BY_M6
  `define AXI_NV_S14_BY_M6 `i_axi_AXI_NV_S14_BY_M6
`endif 

`ifdef i_axi_AXI_NV_S14_BY_M7
  `define AXI_NV_S14_BY_M7 `i_axi_AXI_NV_S14_BY_M7
`endif 

`ifdef i_axi_AXI_NV_S14_BY_M8
  `define AXI_NV_S14_BY_M8 `i_axi_AXI_NV_S14_BY_M8
`endif 

`ifdef i_axi_AXI_NV_S14_BY_M9
  `define AXI_NV_S14_BY_M9 `i_axi_AXI_NV_S14_BY_M9
`endif 

`ifdef i_axi_AXI_NV_S14_BY_M10
  `define AXI_NV_S14_BY_M10 `i_axi_AXI_NV_S14_BY_M10
`endif 

`ifdef i_axi_AXI_NV_S14_BY_M11
  `define AXI_NV_S14_BY_M11 `i_axi_AXI_NV_S14_BY_M11
`endif 

`ifdef i_axi_AXI_NV_S14_BY_M12
  `define AXI_NV_S14_BY_M12 `i_axi_AXI_NV_S14_BY_M12
`endif 

`ifdef i_axi_AXI_NV_S14_BY_M13
  `define AXI_NV_S14_BY_M13 `i_axi_AXI_NV_S14_BY_M13
`endif 

`ifdef i_axi_AXI_NV_S14_BY_M14
  `define AXI_NV_S14_BY_M14 `i_axi_AXI_NV_S14_BY_M14
`endif 

`ifdef i_axi_AXI_NV_S14_BY_M15
  `define AXI_NV_S14_BY_M15 `i_axi_AXI_NV_S14_BY_M15
`endif 

`ifdef i_axi_AXI_NV_S14_BY_M16
  `define AXI_NV_S14_BY_M16 `i_axi_AXI_NV_S14_BY_M16
`endif 

`ifdef i_axi_AXI_NV_S15_BY_M1
  `define AXI_NV_S15_BY_M1 `i_axi_AXI_NV_S15_BY_M1
`endif 

`ifdef i_axi_AXI_NV_S15_BY_M2
  `define AXI_NV_S15_BY_M2 `i_axi_AXI_NV_S15_BY_M2
`endif 

`ifdef i_axi_AXI_NV_S15_BY_M3
  `define AXI_NV_S15_BY_M3 `i_axi_AXI_NV_S15_BY_M3
`endif 

`ifdef i_axi_AXI_NV_S15_BY_M4
  `define AXI_NV_S15_BY_M4 `i_axi_AXI_NV_S15_BY_M4
`endif 

`ifdef i_axi_AXI_NV_S15_BY_M5
  `define AXI_NV_S15_BY_M5 `i_axi_AXI_NV_S15_BY_M5
`endif 

`ifdef i_axi_AXI_NV_S15_BY_M6
  `define AXI_NV_S15_BY_M6 `i_axi_AXI_NV_S15_BY_M6
`endif 

`ifdef i_axi_AXI_NV_S15_BY_M7
  `define AXI_NV_S15_BY_M7 `i_axi_AXI_NV_S15_BY_M7
`endif 

`ifdef i_axi_AXI_NV_S15_BY_M8
  `define AXI_NV_S15_BY_M8 `i_axi_AXI_NV_S15_BY_M8
`endif 

`ifdef i_axi_AXI_NV_S15_BY_M9
  `define AXI_NV_S15_BY_M9 `i_axi_AXI_NV_S15_BY_M9
`endif 

`ifdef i_axi_AXI_NV_S15_BY_M10
  `define AXI_NV_S15_BY_M10 `i_axi_AXI_NV_S15_BY_M10
`endif 

`ifdef i_axi_AXI_NV_S15_BY_M11
  `define AXI_NV_S15_BY_M11 `i_axi_AXI_NV_S15_BY_M11
`endif 

`ifdef i_axi_AXI_NV_S15_BY_M12
  `define AXI_NV_S15_BY_M12 `i_axi_AXI_NV_S15_BY_M12
`endif 

`ifdef i_axi_AXI_NV_S15_BY_M13
  `define AXI_NV_S15_BY_M13 `i_axi_AXI_NV_S15_BY_M13
`endif 

`ifdef i_axi_AXI_NV_S15_BY_M14
  `define AXI_NV_S15_BY_M14 `i_axi_AXI_NV_S15_BY_M14
`endif 

`ifdef i_axi_AXI_NV_S15_BY_M15
  `define AXI_NV_S15_BY_M15 `i_axi_AXI_NV_S15_BY_M15
`endif 

`ifdef i_axi_AXI_NV_S15_BY_M16
  `define AXI_NV_S15_BY_M16 `i_axi_AXI_NV_S15_BY_M16
`endif 

`ifdef i_axi_AXI_NV_S16_BY_M1
  `define AXI_NV_S16_BY_M1 `i_axi_AXI_NV_S16_BY_M1
`endif 

`ifdef i_axi_AXI_NV_S16_BY_M2
  `define AXI_NV_S16_BY_M2 `i_axi_AXI_NV_S16_BY_M2
`endif 

`ifdef i_axi_AXI_NV_S16_BY_M3
  `define AXI_NV_S16_BY_M3 `i_axi_AXI_NV_S16_BY_M3
`endif 

`ifdef i_axi_AXI_NV_S16_BY_M4
  `define AXI_NV_S16_BY_M4 `i_axi_AXI_NV_S16_BY_M4
`endif 

`ifdef i_axi_AXI_NV_S16_BY_M5
  `define AXI_NV_S16_BY_M5 `i_axi_AXI_NV_S16_BY_M5
`endif 

`ifdef i_axi_AXI_NV_S16_BY_M6
  `define AXI_NV_S16_BY_M6 `i_axi_AXI_NV_S16_BY_M6
`endif 

`ifdef i_axi_AXI_NV_S16_BY_M7
  `define AXI_NV_S16_BY_M7 `i_axi_AXI_NV_S16_BY_M7
`endif 

`ifdef i_axi_AXI_NV_S16_BY_M8
  `define AXI_NV_S16_BY_M8 `i_axi_AXI_NV_S16_BY_M8
`endif 

`ifdef i_axi_AXI_NV_S16_BY_M9
  `define AXI_NV_S16_BY_M9 `i_axi_AXI_NV_S16_BY_M9
`endif 

`ifdef i_axi_AXI_NV_S16_BY_M10
  `define AXI_NV_S16_BY_M10 `i_axi_AXI_NV_S16_BY_M10
`endif 

`ifdef i_axi_AXI_NV_S16_BY_M11
  `define AXI_NV_S16_BY_M11 `i_axi_AXI_NV_S16_BY_M11
`endif 

`ifdef i_axi_AXI_NV_S16_BY_M12
  `define AXI_NV_S16_BY_M12 `i_axi_AXI_NV_S16_BY_M12
`endif 

`ifdef i_axi_AXI_NV_S16_BY_M13
  `define AXI_NV_S16_BY_M13 `i_axi_AXI_NV_S16_BY_M13
`endif 

`ifdef i_axi_AXI_NV_S16_BY_M14
  `define AXI_NV_S16_BY_M14 `i_axi_AXI_NV_S16_BY_M14
`endif 

`ifdef i_axi_AXI_NV_S16_BY_M15
  `define AXI_NV_S16_BY_M15 `i_axi_AXI_NV_S16_BY_M15
`endif 

`ifdef i_axi_AXI_NV_S16_BY_M16
  `define AXI_NV_S16_BY_M16 `i_axi_AXI_NV_S16_BY_M16
`endif 

`ifdef i_axi_AXI_NV_S1_BY_ANY_M
  `define AXI_NV_S1_BY_ANY_M `i_axi_AXI_NV_S1_BY_ANY_M
`endif 

`ifdef i_axi_AXI_NV_S2_BY_ANY_M
  `define AXI_NV_S2_BY_ANY_M `i_axi_AXI_NV_S2_BY_ANY_M
`endif 

`ifdef i_axi_AXI_NV_S3_BY_ANY_M
  `define AXI_NV_S3_BY_ANY_M `i_axi_AXI_NV_S3_BY_ANY_M
`endif 

`ifdef i_axi_AXI_NV_S4_BY_ANY_M
  `define AXI_NV_S4_BY_ANY_M `i_axi_AXI_NV_S4_BY_ANY_M
`endif 

`ifdef i_axi_AXI_NV_S5_BY_ANY_M
  `define AXI_NV_S5_BY_ANY_M `i_axi_AXI_NV_S5_BY_ANY_M
`endif 

`ifdef i_axi_AXI_NV_S6_BY_ANY_M
  `define AXI_NV_S6_BY_ANY_M `i_axi_AXI_NV_S6_BY_ANY_M
`endif 

`ifdef i_axi_AXI_NV_S7_BY_ANY_M
  `define AXI_NV_S7_BY_ANY_M `i_axi_AXI_NV_S7_BY_ANY_M
`endif 

`ifdef i_axi_AXI_NV_S8_BY_ANY_M
  `define AXI_NV_S8_BY_ANY_M `i_axi_AXI_NV_S8_BY_ANY_M
`endif 

`ifdef i_axi_AXI_NV_S9_BY_ANY_M
  `define AXI_NV_S9_BY_ANY_M `i_axi_AXI_NV_S9_BY_ANY_M
`endif 

`ifdef i_axi_AXI_NV_S10_BY_ANY_M
  `define AXI_NV_S10_BY_ANY_M `i_axi_AXI_NV_S10_BY_ANY_M
`endif 

`ifdef i_axi_AXI_NV_S11_BY_ANY_M
  `define AXI_NV_S11_BY_ANY_M `i_axi_AXI_NV_S11_BY_ANY_M
`endif 

`ifdef i_axi_AXI_NV_S12_BY_ANY_M
  `define AXI_NV_S12_BY_ANY_M `i_axi_AXI_NV_S12_BY_ANY_M
`endif 

`ifdef i_axi_AXI_NV_S13_BY_ANY_M
  `define AXI_NV_S13_BY_ANY_M `i_axi_AXI_NV_S13_BY_ANY_M
`endif 

`ifdef i_axi_AXI_NV_S14_BY_ANY_M
  `define AXI_NV_S14_BY_ANY_M `i_axi_AXI_NV_S14_BY_ANY_M
`endif 

`ifdef i_axi_AXI_NV_S15_BY_ANY_M
  `define AXI_NV_S15_BY_ANY_M `i_axi_AXI_NV_S15_BY_ANY_M
`endif 

`ifdef i_axi_AXI_NV_S16_BY_ANY_M
  `define AXI_NV_S16_BY_ANY_M `i_axi_AXI_NV_S16_BY_ANY_M
`endif 

`ifdef i_axi_AXI_BV_S0_BY_M1
  `define AXI_BV_S0_BY_M1 `i_axi_AXI_BV_S0_BY_M1
`endif 

`ifdef i_axi_AXI_BV_S0_BY_M2
  `define AXI_BV_S0_BY_M2 `i_axi_AXI_BV_S0_BY_M2
`endif 

`ifdef i_axi_AXI_BV_S0_BY_M3
  `define AXI_BV_S0_BY_M3 `i_axi_AXI_BV_S0_BY_M3
`endif 

`ifdef i_axi_AXI_BV_S0_BY_M4
  `define AXI_BV_S0_BY_M4 `i_axi_AXI_BV_S0_BY_M4
`endif 

`ifdef i_axi_AXI_BV_S0_BY_M5
  `define AXI_BV_S0_BY_M5 `i_axi_AXI_BV_S0_BY_M5
`endif 

`ifdef i_axi_AXI_BV_S0_BY_M6
  `define AXI_BV_S0_BY_M6 `i_axi_AXI_BV_S0_BY_M6
`endif 

`ifdef i_axi_AXI_BV_S0_BY_M7
  `define AXI_BV_S0_BY_M7 `i_axi_AXI_BV_S0_BY_M7
`endif 

`ifdef i_axi_AXI_BV_S0_BY_M8
  `define AXI_BV_S0_BY_M8 `i_axi_AXI_BV_S0_BY_M8
`endif 

`ifdef i_axi_AXI_BV_S0_BY_M9
  `define AXI_BV_S0_BY_M9 `i_axi_AXI_BV_S0_BY_M9
`endif 

`ifdef i_axi_AXI_BV_S0_BY_M10
  `define AXI_BV_S0_BY_M10 `i_axi_AXI_BV_S0_BY_M10
`endif 

`ifdef i_axi_AXI_BV_S0_BY_M11
  `define AXI_BV_S0_BY_M11 `i_axi_AXI_BV_S0_BY_M11
`endif 

`ifdef i_axi_AXI_BV_S0_BY_M12
  `define AXI_BV_S0_BY_M12 `i_axi_AXI_BV_S0_BY_M12
`endif 

`ifdef i_axi_AXI_BV_S0_BY_M13
  `define AXI_BV_S0_BY_M13 `i_axi_AXI_BV_S0_BY_M13
`endif 

`ifdef i_axi_AXI_BV_S0_BY_M14
  `define AXI_BV_S0_BY_M14 `i_axi_AXI_BV_S0_BY_M14
`endif 

`ifdef i_axi_AXI_BV_S0_BY_M15
  `define AXI_BV_S0_BY_M15 `i_axi_AXI_BV_S0_BY_M15
`endif 

`ifdef i_axi_AXI_BV_S0_BY_M16
  `define AXI_BV_S0_BY_M16 `i_axi_AXI_BV_S0_BY_M16
`endif 

`ifdef i_axi_AXI_BV_S1_BY_M1
  `define AXI_BV_S1_BY_M1 `i_axi_AXI_BV_S1_BY_M1
`endif 

`ifdef i_axi_AXI_BV_S1_BY_M2
  `define AXI_BV_S1_BY_M2 `i_axi_AXI_BV_S1_BY_M2
`endif 

`ifdef i_axi_AXI_BV_S1_BY_M3
  `define AXI_BV_S1_BY_M3 `i_axi_AXI_BV_S1_BY_M3
`endif 

`ifdef i_axi_AXI_BV_S1_BY_M4
  `define AXI_BV_S1_BY_M4 `i_axi_AXI_BV_S1_BY_M4
`endif 

`ifdef i_axi_AXI_BV_S1_BY_M5
  `define AXI_BV_S1_BY_M5 `i_axi_AXI_BV_S1_BY_M5
`endif 

`ifdef i_axi_AXI_BV_S1_BY_M6
  `define AXI_BV_S1_BY_M6 `i_axi_AXI_BV_S1_BY_M6
`endif 

`ifdef i_axi_AXI_BV_S1_BY_M7
  `define AXI_BV_S1_BY_M7 `i_axi_AXI_BV_S1_BY_M7
`endif 

`ifdef i_axi_AXI_BV_S1_BY_M8
  `define AXI_BV_S1_BY_M8 `i_axi_AXI_BV_S1_BY_M8
`endif 

`ifdef i_axi_AXI_BV_S1_BY_M9
  `define AXI_BV_S1_BY_M9 `i_axi_AXI_BV_S1_BY_M9
`endif 

`ifdef i_axi_AXI_BV_S1_BY_M10
  `define AXI_BV_S1_BY_M10 `i_axi_AXI_BV_S1_BY_M10
`endif 

`ifdef i_axi_AXI_BV_S1_BY_M11
  `define AXI_BV_S1_BY_M11 `i_axi_AXI_BV_S1_BY_M11
`endif 

`ifdef i_axi_AXI_BV_S1_BY_M12
  `define AXI_BV_S1_BY_M12 `i_axi_AXI_BV_S1_BY_M12
`endif 

`ifdef i_axi_AXI_BV_S1_BY_M13
  `define AXI_BV_S1_BY_M13 `i_axi_AXI_BV_S1_BY_M13
`endif 

`ifdef i_axi_AXI_BV_S1_BY_M14
  `define AXI_BV_S1_BY_M14 `i_axi_AXI_BV_S1_BY_M14
`endif 

`ifdef i_axi_AXI_BV_S1_BY_M15
  `define AXI_BV_S1_BY_M15 `i_axi_AXI_BV_S1_BY_M15
`endif 

`ifdef i_axi_AXI_BV_S1_BY_M16
  `define AXI_BV_S1_BY_M16 `i_axi_AXI_BV_S1_BY_M16
`endif 

`ifdef i_axi_AXI_BV_S2_BY_M1
  `define AXI_BV_S2_BY_M1 `i_axi_AXI_BV_S2_BY_M1
`endif 

`ifdef i_axi_AXI_BV_S2_BY_M2
  `define AXI_BV_S2_BY_M2 `i_axi_AXI_BV_S2_BY_M2
`endif 

`ifdef i_axi_AXI_BV_S2_BY_M3
  `define AXI_BV_S2_BY_M3 `i_axi_AXI_BV_S2_BY_M3
`endif 

`ifdef i_axi_AXI_BV_S2_BY_M4
  `define AXI_BV_S2_BY_M4 `i_axi_AXI_BV_S2_BY_M4
`endif 

`ifdef i_axi_AXI_BV_S2_BY_M5
  `define AXI_BV_S2_BY_M5 `i_axi_AXI_BV_S2_BY_M5
`endif 

`ifdef i_axi_AXI_BV_S2_BY_M6
  `define AXI_BV_S2_BY_M6 `i_axi_AXI_BV_S2_BY_M6
`endif 

`ifdef i_axi_AXI_BV_S2_BY_M7
  `define AXI_BV_S2_BY_M7 `i_axi_AXI_BV_S2_BY_M7
`endif 

`ifdef i_axi_AXI_BV_S2_BY_M8
  `define AXI_BV_S2_BY_M8 `i_axi_AXI_BV_S2_BY_M8
`endif 

`ifdef i_axi_AXI_BV_S2_BY_M9
  `define AXI_BV_S2_BY_M9 `i_axi_AXI_BV_S2_BY_M9
`endif 

`ifdef i_axi_AXI_BV_S2_BY_M10
  `define AXI_BV_S2_BY_M10 `i_axi_AXI_BV_S2_BY_M10
`endif 

`ifdef i_axi_AXI_BV_S2_BY_M11
  `define AXI_BV_S2_BY_M11 `i_axi_AXI_BV_S2_BY_M11
`endif 

`ifdef i_axi_AXI_BV_S2_BY_M12
  `define AXI_BV_S2_BY_M12 `i_axi_AXI_BV_S2_BY_M12
`endif 

`ifdef i_axi_AXI_BV_S2_BY_M13
  `define AXI_BV_S2_BY_M13 `i_axi_AXI_BV_S2_BY_M13
`endif 

`ifdef i_axi_AXI_BV_S2_BY_M14
  `define AXI_BV_S2_BY_M14 `i_axi_AXI_BV_S2_BY_M14
`endif 

`ifdef i_axi_AXI_BV_S2_BY_M15
  `define AXI_BV_S2_BY_M15 `i_axi_AXI_BV_S2_BY_M15
`endif 

`ifdef i_axi_AXI_BV_S2_BY_M16
  `define AXI_BV_S2_BY_M16 `i_axi_AXI_BV_S2_BY_M16
`endif 

`ifdef i_axi_AXI_BV_S3_BY_M1
  `define AXI_BV_S3_BY_M1 `i_axi_AXI_BV_S3_BY_M1
`endif 

`ifdef i_axi_AXI_BV_S3_BY_M2
  `define AXI_BV_S3_BY_M2 `i_axi_AXI_BV_S3_BY_M2
`endif 

`ifdef i_axi_AXI_BV_S3_BY_M3
  `define AXI_BV_S3_BY_M3 `i_axi_AXI_BV_S3_BY_M3
`endif 

`ifdef i_axi_AXI_BV_S3_BY_M4
  `define AXI_BV_S3_BY_M4 `i_axi_AXI_BV_S3_BY_M4
`endif 

`ifdef i_axi_AXI_BV_S3_BY_M5
  `define AXI_BV_S3_BY_M5 `i_axi_AXI_BV_S3_BY_M5
`endif 

`ifdef i_axi_AXI_BV_S3_BY_M6
  `define AXI_BV_S3_BY_M6 `i_axi_AXI_BV_S3_BY_M6
`endif 

`ifdef i_axi_AXI_BV_S3_BY_M7
  `define AXI_BV_S3_BY_M7 `i_axi_AXI_BV_S3_BY_M7
`endif 

`ifdef i_axi_AXI_BV_S3_BY_M8
  `define AXI_BV_S3_BY_M8 `i_axi_AXI_BV_S3_BY_M8
`endif 

`ifdef i_axi_AXI_BV_S3_BY_M9
  `define AXI_BV_S3_BY_M9 `i_axi_AXI_BV_S3_BY_M9
`endif 

`ifdef i_axi_AXI_BV_S3_BY_M10
  `define AXI_BV_S3_BY_M10 `i_axi_AXI_BV_S3_BY_M10
`endif 

`ifdef i_axi_AXI_BV_S3_BY_M11
  `define AXI_BV_S3_BY_M11 `i_axi_AXI_BV_S3_BY_M11
`endif 

`ifdef i_axi_AXI_BV_S3_BY_M12
  `define AXI_BV_S3_BY_M12 `i_axi_AXI_BV_S3_BY_M12
`endif 

`ifdef i_axi_AXI_BV_S3_BY_M13
  `define AXI_BV_S3_BY_M13 `i_axi_AXI_BV_S3_BY_M13
`endif 

`ifdef i_axi_AXI_BV_S3_BY_M14
  `define AXI_BV_S3_BY_M14 `i_axi_AXI_BV_S3_BY_M14
`endif 

`ifdef i_axi_AXI_BV_S3_BY_M15
  `define AXI_BV_S3_BY_M15 `i_axi_AXI_BV_S3_BY_M15
`endif 

`ifdef i_axi_AXI_BV_S3_BY_M16
  `define AXI_BV_S3_BY_M16 `i_axi_AXI_BV_S3_BY_M16
`endif 

`ifdef i_axi_AXI_BV_S4_BY_M1
  `define AXI_BV_S4_BY_M1 `i_axi_AXI_BV_S4_BY_M1
`endif 

`ifdef i_axi_AXI_BV_S4_BY_M2
  `define AXI_BV_S4_BY_M2 `i_axi_AXI_BV_S4_BY_M2
`endif 

`ifdef i_axi_AXI_BV_S4_BY_M3
  `define AXI_BV_S4_BY_M3 `i_axi_AXI_BV_S4_BY_M3
`endif 

`ifdef i_axi_AXI_BV_S4_BY_M4
  `define AXI_BV_S4_BY_M4 `i_axi_AXI_BV_S4_BY_M4
`endif 

`ifdef i_axi_AXI_BV_S4_BY_M5
  `define AXI_BV_S4_BY_M5 `i_axi_AXI_BV_S4_BY_M5
`endif 

`ifdef i_axi_AXI_BV_S4_BY_M6
  `define AXI_BV_S4_BY_M6 `i_axi_AXI_BV_S4_BY_M6
`endif 

`ifdef i_axi_AXI_BV_S4_BY_M7
  `define AXI_BV_S4_BY_M7 `i_axi_AXI_BV_S4_BY_M7
`endif 

`ifdef i_axi_AXI_BV_S4_BY_M8
  `define AXI_BV_S4_BY_M8 `i_axi_AXI_BV_S4_BY_M8
`endif 

`ifdef i_axi_AXI_BV_S4_BY_M9
  `define AXI_BV_S4_BY_M9 `i_axi_AXI_BV_S4_BY_M9
`endif 

`ifdef i_axi_AXI_BV_S4_BY_M10
  `define AXI_BV_S4_BY_M10 `i_axi_AXI_BV_S4_BY_M10
`endif 

`ifdef i_axi_AXI_BV_S4_BY_M11
  `define AXI_BV_S4_BY_M11 `i_axi_AXI_BV_S4_BY_M11
`endif 

`ifdef i_axi_AXI_BV_S4_BY_M12
  `define AXI_BV_S4_BY_M12 `i_axi_AXI_BV_S4_BY_M12
`endif 

`ifdef i_axi_AXI_BV_S4_BY_M13
  `define AXI_BV_S4_BY_M13 `i_axi_AXI_BV_S4_BY_M13
`endif 

`ifdef i_axi_AXI_BV_S4_BY_M14
  `define AXI_BV_S4_BY_M14 `i_axi_AXI_BV_S4_BY_M14
`endif 

`ifdef i_axi_AXI_BV_S4_BY_M15
  `define AXI_BV_S4_BY_M15 `i_axi_AXI_BV_S4_BY_M15
`endif 

`ifdef i_axi_AXI_BV_S4_BY_M16
  `define AXI_BV_S4_BY_M16 `i_axi_AXI_BV_S4_BY_M16
`endif 

`ifdef i_axi_AXI_BV_S5_BY_M1
  `define AXI_BV_S5_BY_M1 `i_axi_AXI_BV_S5_BY_M1
`endif 

`ifdef i_axi_AXI_BV_S5_BY_M2
  `define AXI_BV_S5_BY_M2 `i_axi_AXI_BV_S5_BY_M2
`endif 

`ifdef i_axi_AXI_BV_S5_BY_M3
  `define AXI_BV_S5_BY_M3 `i_axi_AXI_BV_S5_BY_M3
`endif 

`ifdef i_axi_AXI_BV_S5_BY_M4
  `define AXI_BV_S5_BY_M4 `i_axi_AXI_BV_S5_BY_M4
`endif 

`ifdef i_axi_AXI_BV_S5_BY_M5
  `define AXI_BV_S5_BY_M5 `i_axi_AXI_BV_S5_BY_M5
`endif 

`ifdef i_axi_AXI_BV_S5_BY_M6
  `define AXI_BV_S5_BY_M6 `i_axi_AXI_BV_S5_BY_M6
`endif 

`ifdef i_axi_AXI_BV_S5_BY_M7
  `define AXI_BV_S5_BY_M7 `i_axi_AXI_BV_S5_BY_M7
`endif 

`ifdef i_axi_AXI_BV_S5_BY_M8
  `define AXI_BV_S5_BY_M8 `i_axi_AXI_BV_S5_BY_M8
`endif 

`ifdef i_axi_AXI_BV_S5_BY_M9
  `define AXI_BV_S5_BY_M9 `i_axi_AXI_BV_S5_BY_M9
`endif 

`ifdef i_axi_AXI_BV_S5_BY_M10
  `define AXI_BV_S5_BY_M10 `i_axi_AXI_BV_S5_BY_M10
`endif 

`ifdef i_axi_AXI_BV_S5_BY_M11
  `define AXI_BV_S5_BY_M11 `i_axi_AXI_BV_S5_BY_M11
`endif 

`ifdef i_axi_AXI_BV_S5_BY_M12
  `define AXI_BV_S5_BY_M12 `i_axi_AXI_BV_S5_BY_M12
`endif 

`ifdef i_axi_AXI_BV_S5_BY_M13
  `define AXI_BV_S5_BY_M13 `i_axi_AXI_BV_S5_BY_M13
`endif 

`ifdef i_axi_AXI_BV_S5_BY_M14
  `define AXI_BV_S5_BY_M14 `i_axi_AXI_BV_S5_BY_M14
`endif 

`ifdef i_axi_AXI_BV_S5_BY_M15
  `define AXI_BV_S5_BY_M15 `i_axi_AXI_BV_S5_BY_M15
`endif 

`ifdef i_axi_AXI_BV_S5_BY_M16
  `define AXI_BV_S5_BY_M16 `i_axi_AXI_BV_S5_BY_M16
`endif 

`ifdef i_axi_AXI_BV_S6_BY_M1
  `define AXI_BV_S6_BY_M1 `i_axi_AXI_BV_S6_BY_M1
`endif 

`ifdef i_axi_AXI_BV_S6_BY_M2
  `define AXI_BV_S6_BY_M2 `i_axi_AXI_BV_S6_BY_M2
`endif 

`ifdef i_axi_AXI_BV_S6_BY_M3
  `define AXI_BV_S6_BY_M3 `i_axi_AXI_BV_S6_BY_M3
`endif 

`ifdef i_axi_AXI_BV_S6_BY_M4
  `define AXI_BV_S6_BY_M4 `i_axi_AXI_BV_S6_BY_M4
`endif 

`ifdef i_axi_AXI_BV_S6_BY_M5
  `define AXI_BV_S6_BY_M5 `i_axi_AXI_BV_S6_BY_M5
`endif 

`ifdef i_axi_AXI_BV_S6_BY_M6
  `define AXI_BV_S6_BY_M6 `i_axi_AXI_BV_S6_BY_M6
`endif 

`ifdef i_axi_AXI_BV_S6_BY_M7
  `define AXI_BV_S6_BY_M7 `i_axi_AXI_BV_S6_BY_M7
`endif 

`ifdef i_axi_AXI_BV_S6_BY_M8
  `define AXI_BV_S6_BY_M8 `i_axi_AXI_BV_S6_BY_M8
`endif 

`ifdef i_axi_AXI_BV_S6_BY_M9
  `define AXI_BV_S6_BY_M9 `i_axi_AXI_BV_S6_BY_M9
`endif 

`ifdef i_axi_AXI_BV_S6_BY_M10
  `define AXI_BV_S6_BY_M10 `i_axi_AXI_BV_S6_BY_M10
`endif 

`ifdef i_axi_AXI_BV_S6_BY_M11
  `define AXI_BV_S6_BY_M11 `i_axi_AXI_BV_S6_BY_M11
`endif 

`ifdef i_axi_AXI_BV_S6_BY_M12
  `define AXI_BV_S6_BY_M12 `i_axi_AXI_BV_S6_BY_M12
`endif 

`ifdef i_axi_AXI_BV_S6_BY_M13
  `define AXI_BV_S6_BY_M13 `i_axi_AXI_BV_S6_BY_M13
`endif 

`ifdef i_axi_AXI_BV_S6_BY_M14
  `define AXI_BV_S6_BY_M14 `i_axi_AXI_BV_S6_BY_M14
`endif 

`ifdef i_axi_AXI_BV_S6_BY_M15
  `define AXI_BV_S6_BY_M15 `i_axi_AXI_BV_S6_BY_M15
`endif 

`ifdef i_axi_AXI_BV_S6_BY_M16
  `define AXI_BV_S6_BY_M16 `i_axi_AXI_BV_S6_BY_M16
`endif 

`ifdef i_axi_AXI_BV_S7_BY_M1
  `define AXI_BV_S7_BY_M1 `i_axi_AXI_BV_S7_BY_M1
`endif 

`ifdef i_axi_AXI_BV_S7_BY_M2
  `define AXI_BV_S7_BY_M2 `i_axi_AXI_BV_S7_BY_M2
`endif 

`ifdef i_axi_AXI_BV_S7_BY_M3
  `define AXI_BV_S7_BY_M3 `i_axi_AXI_BV_S7_BY_M3
`endif 

`ifdef i_axi_AXI_BV_S7_BY_M4
  `define AXI_BV_S7_BY_M4 `i_axi_AXI_BV_S7_BY_M4
`endif 

`ifdef i_axi_AXI_BV_S7_BY_M5
  `define AXI_BV_S7_BY_M5 `i_axi_AXI_BV_S7_BY_M5
`endif 

`ifdef i_axi_AXI_BV_S7_BY_M6
  `define AXI_BV_S7_BY_M6 `i_axi_AXI_BV_S7_BY_M6
`endif 

`ifdef i_axi_AXI_BV_S7_BY_M7
  `define AXI_BV_S7_BY_M7 `i_axi_AXI_BV_S7_BY_M7
`endif 

`ifdef i_axi_AXI_BV_S7_BY_M8
  `define AXI_BV_S7_BY_M8 `i_axi_AXI_BV_S7_BY_M8
`endif 

`ifdef i_axi_AXI_BV_S7_BY_M9
  `define AXI_BV_S7_BY_M9 `i_axi_AXI_BV_S7_BY_M9
`endif 

`ifdef i_axi_AXI_BV_S7_BY_M10
  `define AXI_BV_S7_BY_M10 `i_axi_AXI_BV_S7_BY_M10
`endif 

`ifdef i_axi_AXI_BV_S7_BY_M11
  `define AXI_BV_S7_BY_M11 `i_axi_AXI_BV_S7_BY_M11
`endif 

`ifdef i_axi_AXI_BV_S7_BY_M12
  `define AXI_BV_S7_BY_M12 `i_axi_AXI_BV_S7_BY_M12
`endif 

`ifdef i_axi_AXI_BV_S7_BY_M13
  `define AXI_BV_S7_BY_M13 `i_axi_AXI_BV_S7_BY_M13
`endif 

`ifdef i_axi_AXI_BV_S7_BY_M14
  `define AXI_BV_S7_BY_M14 `i_axi_AXI_BV_S7_BY_M14
`endif 

`ifdef i_axi_AXI_BV_S7_BY_M15
  `define AXI_BV_S7_BY_M15 `i_axi_AXI_BV_S7_BY_M15
`endif 

`ifdef i_axi_AXI_BV_S7_BY_M16
  `define AXI_BV_S7_BY_M16 `i_axi_AXI_BV_S7_BY_M16
`endif 

`ifdef i_axi_AXI_BV_S8_BY_M1
  `define AXI_BV_S8_BY_M1 `i_axi_AXI_BV_S8_BY_M1
`endif 

`ifdef i_axi_AXI_BV_S8_BY_M2
  `define AXI_BV_S8_BY_M2 `i_axi_AXI_BV_S8_BY_M2
`endif 

`ifdef i_axi_AXI_BV_S8_BY_M3
  `define AXI_BV_S8_BY_M3 `i_axi_AXI_BV_S8_BY_M3
`endif 

`ifdef i_axi_AXI_BV_S8_BY_M4
  `define AXI_BV_S8_BY_M4 `i_axi_AXI_BV_S8_BY_M4
`endif 

`ifdef i_axi_AXI_BV_S8_BY_M5
  `define AXI_BV_S8_BY_M5 `i_axi_AXI_BV_S8_BY_M5
`endif 

`ifdef i_axi_AXI_BV_S8_BY_M6
  `define AXI_BV_S8_BY_M6 `i_axi_AXI_BV_S8_BY_M6
`endif 

`ifdef i_axi_AXI_BV_S8_BY_M7
  `define AXI_BV_S8_BY_M7 `i_axi_AXI_BV_S8_BY_M7
`endif 

`ifdef i_axi_AXI_BV_S8_BY_M8
  `define AXI_BV_S8_BY_M8 `i_axi_AXI_BV_S8_BY_M8
`endif 

`ifdef i_axi_AXI_BV_S8_BY_M9
  `define AXI_BV_S8_BY_M9 `i_axi_AXI_BV_S8_BY_M9
`endif 

`ifdef i_axi_AXI_BV_S8_BY_M10
  `define AXI_BV_S8_BY_M10 `i_axi_AXI_BV_S8_BY_M10
`endif 

`ifdef i_axi_AXI_BV_S8_BY_M11
  `define AXI_BV_S8_BY_M11 `i_axi_AXI_BV_S8_BY_M11
`endif 

`ifdef i_axi_AXI_BV_S8_BY_M12
  `define AXI_BV_S8_BY_M12 `i_axi_AXI_BV_S8_BY_M12
`endif 

`ifdef i_axi_AXI_BV_S8_BY_M13
  `define AXI_BV_S8_BY_M13 `i_axi_AXI_BV_S8_BY_M13
`endif 

`ifdef i_axi_AXI_BV_S8_BY_M14
  `define AXI_BV_S8_BY_M14 `i_axi_AXI_BV_S8_BY_M14
`endif 

`ifdef i_axi_AXI_BV_S8_BY_M15
  `define AXI_BV_S8_BY_M15 `i_axi_AXI_BV_S8_BY_M15
`endif 

`ifdef i_axi_AXI_BV_S8_BY_M16
  `define AXI_BV_S8_BY_M16 `i_axi_AXI_BV_S8_BY_M16
`endif 

`ifdef i_axi_AXI_BV_S9_BY_M1
  `define AXI_BV_S9_BY_M1 `i_axi_AXI_BV_S9_BY_M1
`endif 

`ifdef i_axi_AXI_BV_S9_BY_M2
  `define AXI_BV_S9_BY_M2 `i_axi_AXI_BV_S9_BY_M2
`endif 

`ifdef i_axi_AXI_BV_S9_BY_M3
  `define AXI_BV_S9_BY_M3 `i_axi_AXI_BV_S9_BY_M3
`endif 

`ifdef i_axi_AXI_BV_S9_BY_M4
  `define AXI_BV_S9_BY_M4 `i_axi_AXI_BV_S9_BY_M4
`endif 

`ifdef i_axi_AXI_BV_S9_BY_M5
  `define AXI_BV_S9_BY_M5 `i_axi_AXI_BV_S9_BY_M5
`endif 

`ifdef i_axi_AXI_BV_S9_BY_M6
  `define AXI_BV_S9_BY_M6 `i_axi_AXI_BV_S9_BY_M6
`endif 

`ifdef i_axi_AXI_BV_S9_BY_M7
  `define AXI_BV_S9_BY_M7 `i_axi_AXI_BV_S9_BY_M7
`endif 

`ifdef i_axi_AXI_BV_S9_BY_M8
  `define AXI_BV_S9_BY_M8 `i_axi_AXI_BV_S9_BY_M8
`endif 

`ifdef i_axi_AXI_BV_S9_BY_M9
  `define AXI_BV_S9_BY_M9 `i_axi_AXI_BV_S9_BY_M9
`endif 

`ifdef i_axi_AXI_BV_S9_BY_M10
  `define AXI_BV_S9_BY_M10 `i_axi_AXI_BV_S9_BY_M10
`endif 

`ifdef i_axi_AXI_BV_S9_BY_M11
  `define AXI_BV_S9_BY_M11 `i_axi_AXI_BV_S9_BY_M11
`endif 

`ifdef i_axi_AXI_BV_S9_BY_M12
  `define AXI_BV_S9_BY_M12 `i_axi_AXI_BV_S9_BY_M12
`endif 

`ifdef i_axi_AXI_BV_S9_BY_M13
  `define AXI_BV_S9_BY_M13 `i_axi_AXI_BV_S9_BY_M13
`endif 

`ifdef i_axi_AXI_BV_S9_BY_M14
  `define AXI_BV_S9_BY_M14 `i_axi_AXI_BV_S9_BY_M14
`endif 

`ifdef i_axi_AXI_BV_S9_BY_M15
  `define AXI_BV_S9_BY_M15 `i_axi_AXI_BV_S9_BY_M15
`endif 

`ifdef i_axi_AXI_BV_S9_BY_M16
  `define AXI_BV_S9_BY_M16 `i_axi_AXI_BV_S9_BY_M16
`endif 

`ifdef i_axi_AXI_BV_S10_BY_M1
  `define AXI_BV_S10_BY_M1 `i_axi_AXI_BV_S10_BY_M1
`endif 

`ifdef i_axi_AXI_BV_S10_BY_M2
  `define AXI_BV_S10_BY_M2 `i_axi_AXI_BV_S10_BY_M2
`endif 

`ifdef i_axi_AXI_BV_S10_BY_M3
  `define AXI_BV_S10_BY_M3 `i_axi_AXI_BV_S10_BY_M3
`endif 

`ifdef i_axi_AXI_BV_S10_BY_M4
  `define AXI_BV_S10_BY_M4 `i_axi_AXI_BV_S10_BY_M4
`endif 

`ifdef i_axi_AXI_BV_S10_BY_M5
  `define AXI_BV_S10_BY_M5 `i_axi_AXI_BV_S10_BY_M5
`endif 

`ifdef i_axi_AXI_BV_S10_BY_M6
  `define AXI_BV_S10_BY_M6 `i_axi_AXI_BV_S10_BY_M6
`endif 

`ifdef i_axi_AXI_BV_S10_BY_M7
  `define AXI_BV_S10_BY_M7 `i_axi_AXI_BV_S10_BY_M7
`endif 

`ifdef i_axi_AXI_BV_S10_BY_M8
  `define AXI_BV_S10_BY_M8 `i_axi_AXI_BV_S10_BY_M8
`endif 

`ifdef i_axi_AXI_BV_S10_BY_M9
  `define AXI_BV_S10_BY_M9 `i_axi_AXI_BV_S10_BY_M9
`endif 

`ifdef i_axi_AXI_BV_S10_BY_M10
  `define AXI_BV_S10_BY_M10 `i_axi_AXI_BV_S10_BY_M10
`endif 

`ifdef i_axi_AXI_BV_S10_BY_M11
  `define AXI_BV_S10_BY_M11 `i_axi_AXI_BV_S10_BY_M11
`endif 

`ifdef i_axi_AXI_BV_S10_BY_M12
  `define AXI_BV_S10_BY_M12 `i_axi_AXI_BV_S10_BY_M12
`endif 

`ifdef i_axi_AXI_BV_S10_BY_M13
  `define AXI_BV_S10_BY_M13 `i_axi_AXI_BV_S10_BY_M13
`endif 

`ifdef i_axi_AXI_BV_S10_BY_M14
  `define AXI_BV_S10_BY_M14 `i_axi_AXI_BV_S10_BY_M14
`endif 

`ifdef i_axi_AXI_BV_S10_BY_M15
  `define AXI_BV_S10_BY_M15 `i_axi_AXI_BV_S10_BY_M15
`endif 

`ifdef i_axi_AXI_BV_S10_BY_M16
  `define AXI_BV_S10_BY_M16 `i_axi_AXI_BV_S10_BY_M16
`endif 

`ifdef i_axi_AXI_BV_S11_BY_M1
  `define AXI_BV_S11_BY_M1 `i_axi_AXI_BV_S11_BY_M1
`endif 

`ifdef i_axi_AXI_BV_S11_BY_M2
  `define AXI_BV_S11_BY_M2 `i_axi_AXI_BV_S11_BY_M2
`endif 

`ifdef i_axi_AXI_BV_S11_BY_M3
  `define AXI_BV_S11_BY_M3 `i_axi_AXI_BV_S11_BY_M3
`endif 

`ifdef i_axi_AXI_BV_S11_BY_M4
  `define AXI_BV_S11_BY_M4 `i_axi_AXI_BV_S11_BY_M4
`endif 

`ifdef i_axi_AXI_BV_S11_BY_M5
  `define AXI_BV_S11_BY_M5 `i_axi_AXI_BV_S11_BY_M5
`endif 

`ifdef i_axi_AXI_BV_S11_BY_M6
  `define AXI_BV_S11_BY_M6 `i_axi_AXI_BV_S11_BY_M6
`endif 

`ifdef i_axi_AXI_BV_S11_BY_M7
  `define AXI_BV_S11_BY_M7 `i_axi_AXI_BV_S11_BY_M7
`endif 

`ifdef i_axi_AXI_BV_S11_BY_M8
  `define AXI_BV_S11_BY_M8 `i_axi_AXI_BV_S11_BY_M8
`endif 

`ifdef i_axi_AXI_BV_S11_BY_M9
  `define AXI_BV_S11_BY_M9 `i_axi_AXI_BV_S11_BY_M9
`endif 

`ifdef i_axi_AXI_BV_S11_BY_M10
  `define AXI_BV_S11_BY_M10 `i_axi_AXI_BV_S11_BY_M10
`endif 

`ifdef i_axi_AXI_BV_S11_BY_M11
  `define AXI_BV_S11_BY_M11 `i_axi_AXI_BV_S11_BY_M11
`endif 

`ifdef i_axi_AXI_BV_S11_BY_M12
  `define AXI_BV_S11_BY_M12 `i_axi_AXI_BV_S11_BY_M12
`endif 

`ifdef i_axi_AXI_BV_S11_BY_M13
  `define AXI_BV_S11_BY_M13 `i_axi_AXI_BV_S11_BY_M13
`endif 

`ifdef i_axi_AXI_BV_S11_BY_M14
  `define AXI_BV_S11_BY_M14 `i_axi_AXI_BV_S11_BY_M14
`endif 

`ifdef i_axi_AXI_BV_S11_BY_M15
  `define AXI_BV_S11_BY_M15 `i_axi_AXI_BV_S11_BY_M15
`endif 

`ifdef i_axi_AXI_BV_S11_BY_M16
  `define AXI_BV_S11_BY_M16 `i_axi_AXI_BV_S11_BY_M16
`endif 

`ifdef i_axi_AXI_BV_S12_BY_M1
  `define AXI_BV_S12_BY_M1 `i_axi_AXI_BV_S12_BY_M1
`endif 

`ifdef i_axi_AXI_BV_S12_BY_M2
  `define AXI_BV_S12_BY_M2 `i_axi_AXI_BV_S12_BY_M2
`endif 

`ifdef i_axi_AXI_BV_S12_BY_M3
  `define AXI_BV_S12_BY_M3 `i_axi_AXI_BV_S12_BY_M3
`endif 

`ifdef i_axi_AXI_BV_S12_BY_M4
  `define AXI_BV_S12_BY_M4 `i_axi_AXI_BV_S12_BY_M4
`endif 

`ifdef i_axi_AXI_BV_S12_BY_M5
  `define AXI_BV_S12_BY_M5 `i_axi_AXI_BV_S12_BY_M5
`endif 

`ifdef i_axi_AXI_BV_S12_BY_M6
  `define AXI_BV_S12_BY_M6 `i_axi_AXI_BV_S12_BY_M6
`endif 

`ifdef i_axi_AXI_BV_S12_BY_M7
  `define AXI_BV_S12_BY_M7 `i_axi_AXI_BV_S12_BY_M7
`endif 

`ifdef i_axi_AXI_BV_S12_BY_M8
  `define AXI_BV_S12_BY_M8 `i_axi_AXI_BV_S12_BY_M8
`endif 

`ifdef i_axi_AXI_BV_S12_BY_M9
  `define AXI_BV_S12_BY_M9 `i_axi_AXI_BV_S12_BY_M9
`endif 

`ifdef i_axi_AXI_BV_S12_BY_M10
  `define AXI_BV_S12_BY_M10 `i_axi_AXI_BV_S12_BY_M10
`endif 

`ifdef i_axi_AXI_BV_S12_BY_M11
  `define AXI_BV_S12_BY_M11 `i_axi_AXI_BV_S12_BY_M11
`endif 

`ifdef i_axi_AXI_BV_S12_BY_M12
  `define AXI_BV_S12_BY_M12 `i_axi_AXI_BV_S12_BY_M12
`endif 

`ifdef i_axi_AXI_BV_S12_BY_M13
  `define AXI_BV_S12_BY_M13 `i_axi_AXI_BV_S12_BY_M13
`endif 

`ifdef i_axi_AXI_BV_S12_BY_M14
  `define AXI_BV_S12_BY_M14 `i_axi_AXI_BV_S12_BY_M14
`endif 

`ifdef i_axi_AXI_BV_S12_BY_M15
  `define AXI_BV_S12_BY_M15 `i_axi_AXI_BV_S12_BY_M15
`endif 

`ifdef i_axi_AXI_BV_S12_BY_M16
  `define AXI_BV_S12_BY_M16 `i_axi_AXI_BV_S12_BY_M16
`endif 

`ifdef i_axi_AXI_BV_S13_BY_M1
  `define AXI_BV_S13_BY_M1 `i_axi_AXI_BV_S13_BY_M1
`endif 

`ifdef i_axi_AXI_BV_S13_BY_M2
  `define AXI_BV_S13_BY_M2 `i_axi_AXI_BV_S13_BY_M2
`endif 

`ifdef i_axi_AXI_BV_S13_BY_M3
  `define AXI_BV_S13_BY_M3 `i_axi_AXI_BV_S13_BY_M3
`endif 

`ifdef i_axi_AXI_BV_S13_BY_M4
  `define AXI_BV_S13_BY_M4 `i_axi_AXI_BV_S13_BY_M4
`endif 

`ifdef i_axi_AXI_BV_S13_BY_M5
  `define AXI_BV_S13_BY_M5 `i_axi_AXI_BV_S13_BY_M5
`endif 

`ifdef i_axi_AXI_BV_S13_BY_M6
  `define AXI_BV_S13_BY_M6 `i_axi_AXI_BV_S13_BY_M6
`endif 

`ifdef i_axi_AXI_BV_S13_BY_M7
  `define AXI_BV_S13_BY_M7 `i_axi_AXI_BV_S13_BY_M7
`endif 

`ifdef i_axi_AXI_BV_S13_BY_M8
  `define AXI_BV_S13_BY_M8 `i_axi_AXI_BV_S13_BY_M8
`endif 

`ifdef i_axi_AXI_BV_S13_BY_M9
  `define AXI_BV_S13_BY_M9 `i_axi_AXI_BV_S13_BY_M9
`endif 

`ifdef i_axi_AXI_BV_S13_BY_M10
  `define AXI_BV_S13_BY_M10 `i_axi_AXI_BV_S13_BY_M10
`endif 

`ifdef i_axi_AXI_BV_S13_BY_M11
  `define AXI_BV_S13_BY_M11 `i_axi_AXI_BV_S13_BY_M11
`endif 

`ifdef i_axi_AXI_BV_S13_BY_M12
  `define AXI_BV_S13_BY_M12 `i_axi_AXI_BV_S13_BY_M12
`endif 

`ifdef i_axi_AXI_BV_S13_BY_M13
  `define AXI_BV_S13_BY_M13 `i_axi_AXI_BV_S13_BY_M13
`endif 

`ifdef i_axi_AXI_BV_S13_BY_M14
  `define AXI_BV_S13_BY_M14 `i_axi_AXI_BV_S13_BY_M14
`endif 

`ifdef i_axi_AXI_BV_S13_BY_M15
  `define AXI_BV_S13_BY_M15 `i_axi_AXI_BV_S13_BY_M15
`endif 

`ifdef i_axi_AXI_BV_S13_BY_M16
  `define AXI_BV_S13_BY_M16 `i_axi_AXI_BV_S13_BY_M16
`endif 

`ifdef i_axi_AXI_BV_S14_BY_M1
  `define AXI_BV_S14_BY_M1 `i_axi_AXI_BV_S14_BY_M1
`endif 

`ifdef i_axi_AXI_BV_S14_BY_M2
  `define AXI_BV_S14_BY_M2 `i_axi_AXI_BV_S14_BY_M2
`endif 

`ifdef i_axi_AXI_BV_S14_BY_M3
  `define AXI_BV_S14_BY_M3 `i_axi_AXI_BV_S14_BY_M3
`endif 

`ifdef i_axi_AXI_BV_S14_BY_M4
  `define AXI_BV_S14_BY_M4 `i_axi_AXI_BV_S14_BY_M4
`endif 

`ifdef i_axi_AXI_BV_S14_BY_M5
  `define AXI_BV_S14_BY_M5 `i_axi_AXI_BV_S14_BY_M5
`endif 

`ifdef i_axi_AXI_BV_S14_BY_M6
  `define AXI_BV_S14_BY_M6 `i_axi_AXI_BV_S14_BY_M6
`endif 

`ifdef i_axi_AXI_BV_S14_BY_M7
  `define AXI_BV_S14_BY_M7 `i_axi_AXI_BV_S14_BY_M7
`endif 

`ifdef i_axi_AXI_BV_S14_BY_M8
  `define AXI_BV_S14_BY_M8 `i_axi_AXI_BV_S14_BY_M8
`endif 

`ifdef i_axi_AXI_BV_S14_BY_M9
  `define AXI_BV_S14_BY_M9 `i_axi_AXI_BV_S14_BY_M9
`endif 

`ifdef i_axi_AXI_BV_S14_BY_M10
  `define AXI_BV_S14_BY_M10 `i_axi_AXI_BV_S14_BY_M10
`endif 

`ifdef i_axi_AXI_BV_S14_BY_M11
  `define AXI_BV_S14_BY_M11 `i_axi_AXI_BV_S14_BY_M11
`endif 

`ifdef i_axi_AXI_BV_S14_BY_M12
  `define AXI_BV_S14_BY_M12 `i_axi_AXI_BV_S14_BY_M12
`endif 

`ifdef i_axi_AXI_BV_S14_BY_M13
  `define AXI_BV_S14_BY_M13 `i_axi_AXI_BV_S14_BY_M13
`endif 

`ifdef i_axi_AXI_BV_S14_BY_M14
  `define AXI_BV_S14_BY_M14 `i_axi_AXI_BV_S14_BY_M14
`endif 

`ifdef i_axi_AXI_BV_S14_BY_M15
  `define AXI_BV_S14_BY_M15 `i_axi_AXI_BV_S14_BY_M15
`endif 

`ifdef i_axi_AXI_BV_S14_BY_M16
  `define AXI_BV_S14_BY_M16 `i_axi_AXI_BV_S14_BY_M16
`endif 

`ifdef i_axi_AXI_BV_S15_BY_M1
  `define AXI_BV_S15_BY_M1 `i_axi_AXI_BV_S15_BY_M1
`endif 

`ifdef i_axi_AXI_BV_S15_BY_M2
  `define AXI_BV_S15_BY_M2 `i_axi_AXI_BV_S15_BY_M2
`endif 

`ifdef i_axi_AXI_BV_S15_BY_M3
  `define AXI_BV_S15_BY_M3 `i_axi_AXI_BV_S15_BY_M3
`endif 

`ifdef i_axi_AXI_BV_S15_BY_M4
  `define AXI_BV_S15_BY_M4 `i_axi_AXI_BV_S15_BY_M4
`endif 

`ifdef i_axi_AXI_BV_S15_BY_M5
  `define AXI_BV_S15_BY_M5 `i_axi_AXI_BV_S15_BY_M5
`endif 

`ifdef i_axi_AXI_BV_S15_BY_M6
  `define AXI_BV_S15_BY_M6 `i_axi_AXI_BV_S15_BY_M6
`endif 

`ifdef i_axi_AXI_BV_S15_BY_M7
  `define AXI_BV_S15_BY_M7 `i_axi_AXI_BV_S15_BY_M7
`endif 

`ifdef i_axi_AXI_BV_S15_BY_M8
  `define AXI_BV_S15_BY_M8 `i_axi_AXI_BV_S15_BY_M8
`endif 

`ifdef i_axi_AXI_BV_S15_BY_M9
  `define AXI_BV_S15_BY_M9 `i_axi_AXI_BV_S15_BY_M9
`endif 

`ifdef i_axi_AXI_BV_S15_BY_M10
  `define AXI_BV_S15_BY_M10 `i_axi_AXI_BV_S15_BY_M10
`endif 

`ifdef i_axi_AXI_BV_S15_BY_M11
  `define AXI_BV_S15_BY_M11 `i_axi_AXI_BV_S15_BY_M11
`endif 

`ifdef i_axi_AXI_BV_S15_BY_M12
  `define AXI_BV_S15_BY_M12 `i_axi_AXI_BV_S15_BY_M12
`endif 

`ifdef i_axi_AXI_BV_S15_BY_M13
  `define AXI_BV_S15_BY_M13 `i_axi_AXI_BV_S15_BY_M13
`endif 

`ifdef i_axi_AXI_BV_S15_BY_M14
  `define AXI_BV_S15_BY_M14 `i_axi_AXI_BV_S15_BY_M14
`endif 

`ifdef i_axi_AXI_BV_S15_BY_M15
  `define AXI_BV_S15_BY_M15 `i_axi_AXI_BV_S15_BY_M15
`endif 

`ifdef i_axi_AXI_BV_S15_BY_M16
  `define AXI_BV_S15_BY_M16 `i_axi_AXI_BV_S15_BY_M16
`endif 

`ifdef i_axi_AXI_BV_S16_BY_M1
  `define AXI_BV_S16_BY_M1 `i_axi_AXI_BV_S16_BY_M1
`endif 

`ifdef i_axi_AXI_BV_S16_BY_M2
  `define AXI_BV_S16_BY_M2 `i_axi_AXI_BV_S16_BY_M2
`endif 

`ifdef i_axi_AXI_BV_S16_BY_M3
  `define AXI_BV_S16_BY_M3 `i_axi_AXI_BV_S16_BY_M3
`endif 

`ifdef i_axi_AXI_BV_S16_BY_M4
  `define AXI_BV_S16_BY_M4 `i_axi_AXI_BV_S16_BY_M4
`endif 

`ifdef i_axi_AXI_BV_S16_BY_M5
  `define AXI_BV_S16_BY_M5 `i_axi_AXI_BV_S16_BY_M5
`endif 

`ifdef i_axi_AXI_BV_S16_BY_M6
  `define AXI_BV_S16_BY_M6 `i_axi_AXI_BV_S16_BY_M6
`endif 

`ifdef i_axi_AXI_BV_S16_BY_M7
  `define AXI_BV_S16_BY_M7 `i_axi_AXI_BV_S16_BY_M7
`endif 

`ifdef i_axi_AXI_BV_S16_BY_M8
  `define AXI_BV_S16_BY_M8 `i_axi_AXI_BV_S16_BY_M8
`endif 

`ifdef i_axi_AXI_BV_S16_BY_M9
  `define AXI_BV_S16_BY_M9 `i_axi_AXI_BV_S16_BY_M9
`endif 

`ifdef i_axi_AXI_BV_S16_BY_M10
  `define AXI_BV_S16_BY_M10 `i_axi_AXI_BV_S16_BY_M10
`endif 

`ifdef i_axi_AXI_BV_S16_BY_M11
  `define AXI_BV_S16_BY_M11 `i_axi_AXI_BV_S16_BY_M11
`endif 

`ifdef i_axi_AXI_BV_S16_BY_M12
  `define AXI_BV_S16_BY_M12 `i_axi_AXI_BV_S16_BY_M12
`endif 

`ifdef i_axi_AXI_BV_S16_BY_M13
  `define AXI_BV_S16_BY_M13 `i_axi_AXI_BV_S16_BY_M13
`endif 

`ifdef i_axi_AXI_BV_S16_BY_M14
  `define AXI_BV_S16_BY_M14 `i_axi_AXI_BV_S16_BY_M14
`endif 

`ifdef i_axi_AXI_BV_S16_BY_M15
  `define AXI_BV_S16_BY_M15 `i_axi_AXI_BV_S16_BY_M15
`endif 

`ifdef i_axi_AXI_BV_S16_BY_M16
  `define AXI_BV_S16_BY_M16 `i_axi_AXI_BV_S16_BY_M16
`endif 

`ifdef i_axi_AXI_BV_S1_BY_ANY_M
  `define AXI_BV_S1_BY_ANY_M `i_axi_AXI_BV_S1_BY_ANY_M
`endif 

`ifdef i_axi_AXI_BV_S2_BY_ANY_M
  `define AXI_BV_S2_BY_ANY_M `i_axi_AXI_BV_S2_BY_ANY_M
`endif 

`ifdef i_axi_AXI_BV_S3_BY_ANY_M
  `define AXI_BV_S3_BY_ANY_M `i_axi_AXI_BV_S3_BY_ANY_M
`endif 

`ifdef i_axi_AXI_BV_S4_BY_ANY_M
  `define AXI_BV_S4_BY_ANY_M `i_axi_AXI_BV_S4_BY_ANY_M
`endif 

`ifdef i_axi_AXI_BV_S5_BY_ANY_M
  `define AXI_BV_S5_BY_ANY_M `i_axi_AXI_BV_S5_BY_ANY_M
`endif 

`ifdef i_axi_AXI_BV_S6_BY_ANY_M
  `define AXI_BV_S6_BY_ANY_M `i_axi_AXI_BV_S6_BY_ANY_M
`endif 

`ifdef i_axi_AXI_BV_S7_BY_ANY_M
  `define AXI_BV_S7_BY_ANY_M `i_axi_AXI_BV_S7_BY_ANY_M
`endif 

`ifdef i_axi_AXI_BV_S8_BY_ANY_M
  `define AXI_BV_S8_BY_ANY_M `i_axi_AXI_BV_S8_BY_ANY_M
`endif 

`ifdef i_axi_AXI_BV_S9_BY_ANY_M
  `define AXI_BV_S9_BY_ANY_M `i_axi_AXI_BV_S9_BY_ANY_M
`endif 

`ifdef i_axi_AXI_BV_S10_BY_ANY_M
  `define AXI_BV_S10_BY_ANY_M `i_axi_AXI_BV_S10_BY_ANY_M
`endif 

`ifdef i_axi_AXI_BV_S11_BY_ANY_M
  `define AXI_BV_S11_BY_ANY_M `i_axi_AXI_BV_S11_BY_ANY_M
`endif 

`ifdef i_axi_AXI_BV_S12_BY_ANY_M
  `define AXI_BV_S12_BY_ANY_M `i_axi_AXI_BV_S12_BY_ANY_M
`endif 

`ifdef i_axi_AXI_BV_S13_BY_ANY_M
  `define AXI_BV_S13_BY_ANY_M `i_axi_AXI_BV_S13_BY_ANY_M
`endif 

`ifdef i_axi_AXI_BV_S14_BY_ANY_M
  `define AXI_BV_S14_BY_ANY_M `i_axi_AXI_BV_S14_BY_ANY_M
`endif 

`ifdef i_axi_AXI_BV_S15_BY_ANY_M
  `define AXI_BV_S15_BY_ANY_M `i_axi_AXI_BV_S15_BY_ANY_M
`endif 

`ifdef i_axi_AXI_BV_S16_BY_ANY_M
  `define AXI_BV_S16_BY_ANY_M `i_axi_AXI_BV_S16_BY_ANY_M
`endif 

`ifdef i_axi_AXI_VV_S0_BY_M1
  `define AXI_VV_S0_BY_M1 `i_axi_AXI_VV_S0_BY_M1
`endif 

`ifdef i_axi_AXI_V_S0_BY_M1
  `define AXI_V_S0_BY_M1 `i_axi_AXI_V_S0_BY_M1
`endif 

`ifdef i_axi_AXI_VV_S0_BY_M2
  `define AXI_VV_S0_BY_M2 `i_axi_AXI_VV_S0_BY_M2
`endif 

`ifdef i_axi_AXI_V_S0_BY_M2
  `define AXI_V_S0_BY_M2 `i_axi_AXI_V_S0_BY_M2
`endif 

`ifdef i_axi_AXI_VV_S0_BY_M3
  `define AXI_VV_S0_BY_M3 `i_axi_AXI_VV_S0_BY_M3
`endif 

`ifdef i_axi_AXI_VV_S0_BY_M4
  `define AXI_VV_S0_BY_M4 `i_axi_AXI_VV_S0_BY_M4
`endif 

`ifdef i_axi_AXI_VV_S0_BY_M5
  `define AXI_VV_S0_BY_M5 `i_axi_AXI_VV_S0_BY_M5
`endif 

`ifdef i_axi_AXI_VV_S0_BY_M6
  `define AXI_VV_S0_BY_M6 `i_axi_AXI_VV_S0_BY_M6
`endif 

`ifdef i_axi_AXI_VV_S0_BY_M7
  `define AXI_VV_S0_BY_M7 `i_axi_AXI_VV_S0_BY_M7
`endif 

`ifdef i_axi_AXI_VV_S0_BY_M8
  `define AXI_VV_S0_BY_M8 `i_axi_AXI_VV_S0_BY_M8
`endif 

`ifdef i_axi_AXI_VV_S0_BY_M9
  `define AXI_VV_S0_BY_M9 `i_axi_AXI_VV_S0_BY_M9
`endif 

`ifdef i_axi_AXI_VV_S0_BY_M10
  `define AXI_VV_S0_BY_M10 `i_axi_AXI_VV_S0_BY_M10
`endif 

`ifdef i_axi_AXI_VV_S0_BY_M11
  `define AXI_VV_S0_BY_M11 `i_axi_AXI_VV_S0_BY_M11
`endif 

`ifdef i_axi_AXI_VV_S0_BY_M12
  `define AXI_VV_S0_BY_M12 `i_axi_AXI_VV_S0_BY_M12
`endif 

`ifdef i_axi_AXI_VV_S0_BY_M13
  `define AXI_VV_S0_BY_M13 `i_axi_AXI_VV_S0_BY_M13
`endif 

`ifdef i_axi_AXI_VV_S0_BY_M14
  `define AXI_VV_S0_BY_M14 `i_axi_AXI_VV_S0_BY_M14
`endif 

`ifdef i_axi_AXI_VV_S0_BY_M15
  `define AXI_VV_S0_BY_M15 `i_axi_AXI_VV_S0_BY_M15
`endif 

`ifdef i_axi_AXI_VV_S0_BY_M16
  `define AXI_VV_S0_BY_M16 `i_axi_AXI_VV_S0_BY_M16
`endif 

`ifdef i_axi_AXI_VV_S1_BY_M1
  `define AXI_VV_S1_BY_M1 `i_axi_AXI_VV_S1_BY_M1
`endif 

`ifdef i_axi_AXI_V_S1_BY_M1
  `define AXI_V_S1_BY_M1 `i_axi_AXI_V_S1_BY_M1
`endif 

`ifdef i_axi_AXI_VV_S1_BY_M2
  `define AXI_VV_S1_BY_M2 `i_axi_AXI_VV_S1_BY_M2
`endif 

`ifdef i_axi_AXI_V_S1_BY_M2
  `define AXI_V_S1_BY_M2 `i_axi_AXI_V_S1_BY_M2
`endif 

`ifdef i_axi_AXI_VV_S1_BY_M3
  `define AXI_VV_S1_BY_M3 `i_axi_AXI_VV_S1_BY_M3
`endif 

`ifdef i_axi_AXI_VV_S1_BY_M4
  `define AXI_VV_S1_BY_M4 `i_axi_AXI_VV_S1_BY_M4
`endif 

`ifdef i_axi_AXI_VV_S1_BY_M5
  `define AXI_VV_S1_BY_M5 `i_axi_AXI_VV_S1_BY_M5
`endif 

`ifdef i_axi_AXI_VV_S1_BY_M6
  `define AXI_VV_S1_BY_M6 `i_axi_AXI_VV_S1_BY_M6
`endif 

`ifdef i_axi_AXI_VV_S1_BY_M7
  `define AXI_VV_S1_BY_M7 `i_axi_AXI_VV_S1_BY_M7
`endif 

`ifdef i_axi_AXI_VV_S1_BY_M8
  `define AXI_VV_S1_BY_M8 `i_axi_AXI_VV_S1_BY_M8
`endif 

`ifdef i_axi_AXI_VV_S1_BY_M9
  `define AXI_VV_S1_BY_M9 `i_axi_AXI_VV_S1_BY_M9
`endif 

`ifdef i_axi_AXI_VV_S1_BY_M10
  `define AXI_VV_S1_BY_M10 `i_axi_AXI_VV_S1_BY_M10
`endif 

`ifdef i_axi_AXI_VV_S1_BY_M11
  `define AXI_VV_S1_BY_M11 `i_axi_AXI_VV_S1_BY_M11
`endif 

`ifdef i_axi_AXI_VV_S1_BY_M12
  `define AXI_VV_S1_BY_M12 `i_axi_AXI_VV_S1_BY_M12
`endif 

`ifdef i_axi_AXI_VV_S1_BY_M13
  `define AXI_VV_S1_BY_M13 `i_axi_AXI_VV_S1_BY_M13
`endif 

`ifdef i_axi_AXI_VV_S1_BY_M14
  `define AXI_VV_S1_BY_M14 `i_axi_AXI_VV_S1_BY_M14
`endif 

`ifdef i_axi_AXI_VV_S1_BY_M15
  `define AXI_VV_S1_BY_M15 `i_axi_AXI_VV_S1_BY_M15
`endif 

`ifdef i_axi_AXI_VV_S1_BY_M16
  `define AXI_VV_S1_BY_M16 `i_axi_AXI_VV_S1_BY_M16
`endif 

`ifdef i_axi_AXI_VV_S2_BY_M1
  `define AXI_VV_S2_BY_M1 `i_axi_AXI_VV_S2_BY_M1
`endif 

`ifdef i_axi_AXI_V_S2_BY_M1
  `define AXI_V_S2_BY_M1 `i_axi_AXI_V_S2_BY_M1
`endif 

`ifdef i_axi_AXI_VV_S2_BY_M2
  `define AXI_VV_S2_BY_M2 `i_axi_AXI_VV_S2_BY_M2
`endif 

`ifdef i_axi_AXI_V_S2_BY_M2
  `define AXI_V_S2_BY_M2 `i_axi_AXI_V_S2_BY_M2
`endif 

`ifdef i_axi_AXI_VV_S2_BY_M3
  `define AXI_VV_S2_BY_M3 `i_axi_AXI_VV_S2_BY_M3
`endif 

`ifdef i_axi_AXI_VV_S2_BY_M4
  `define AXI_VV_S2_BY_M4 `i_axi_AXI_VV_S2_BY_M4
`endif 

`ifdef i_axi_AXI_VV_S2_BY_M5
  `define AXI_VV_S2_BY_M5 `i_axi_AXI_VV_S2_BY_M5
`endif 

`ifdef i_axi_AXI_VV_S2_BY_M6
  `define AXI_VV_S2_BY_M6 `i_axi_AXI_VV_S2_BY_M6
`endif 

`ifdef i_axi_AXI_VV_S2_BY_M7
  `define AXI_VV_S2_BY_M7 `i_axi_AXI_VV_S2_BY_M7
`endif 

`ifdef i_axi_AXI_VV_S2_BY_M8
  `define AXI_VV_S2_BY_M8 `i_axi_AXI_VV_S2_BY_M8
`endif 

`ifdef i_axi_AXI_VV_S2_BY_M9
  `define AXI_VV_S2_BY_M9 `i_axi_AXI_VV_S2_BY_M9
`endif 

`ifdef i_axi_AXI_VV_S2_BY_M10
  `define AXI_VV_S2_BY_M10 `i_axi_AXI_VV_S2_BY_M10
`endif 

`ifdef i_axi_AXI_VV_S2_BY_M11
  `define AXI_VV_S2_BY_M11 `i_axi_AXI_VV_S2_BY_M11
`endif 

`ifdef i_axi_AXI_VV_S2_BY_M12
  `define AXI_VV_S2_BY_M12 `i_axi_AXI_VV_S2_BY_M12
`endif 

`ifdef i_axi_AXI_VV_S2_BY_M13
  `define AXI_VV_S2_BY_M13 `i_axi_AXI_VV_S2_BY_M13
`endif 

`ifdef i_axi_AXI_VV_S2_BY_M14
  `define AXI_VV_S2_BY_M14 `i_axi_AXI_VV_S2_BY_M14
`endif 

`ifdef i_axi_AXI_VV_S2_BY_M15
  `define AXI_VV_S2_BY_M15 `i_axi_AXI_VV_S2_BY_M15
`endif 

`ifdef i_axi_AXI_VV_S2_BY_M16
  `define AXI_VV_S2_BY_M16 `i_axi_AXI_VV_S2_BY_M16
`endif 

`ifdef i_axi_AXI_VV_S3_BY_M1
  `define AXI_VV_S3_BY_M1 `i_axi_AXI_VV_S3_BY_M1
`endif 

`ifdef i_axi_AXI_V_S3_BY_M1
  `define AXI_V_S3_BY_M1 `i_axi_AXI_V_S3_BY_M1
`endif 

`ifdef i_axi_AXI_VV_S3_BY_M2
  `define AXI_VV_S3_BY_M2 `i_axi_AXI_VV_S3_BY_M2
`endif 

`ifdef i_axi_AXI_V_S3_BY_M2
  `define AXI_V_S3_BY_M2 `i_axi_AXI_V_S3_BY_M2
`endif 

`ifdef i_axi_AXI_VV_S3_BY_M3
  `define AXI_VV_S3_BY_M3 `i_axi_AXI_VV_S3_BY_M3
`endif 

`ifdef i_axi_AXI_VV_S3_BY_M4
  `define AXI_VV_S3_BY_M4 `i_axi_AXI_VV_S3_BY_M4
`endif 

`ifdef i_axi_AXI_VV_S3_BY_M5
  `define AXI_VV_S3_BY_M5 `i_axi_AXI_VV_S3_BY_M5
`endif 

`ifdef i_axi_AXI_VV_S3_BY_M6
  `define AXI_VV_S3_BY_M6 `i_axi_AXI_VV_S3_BY_M6
`endif 

`ifdef i_axi_AXI_VV_S3_BY_M7
  `define AXI_VV_S3_BY_M7 `i_axi_AXI_VV_S3_BY_M7
`endif 

`ifdef i_axi_AXI_VV_S3_BY_M8
  `define AXI_VV_S3_BY_M8 `i_axi_AXI_VV_S3_BY_M8
`endif 

`ifdef i_axi_AXI_VV_S3_BY_M9
  `define AXI_VV_S3_BY_M9 `i_axi_AXI_VV_S3_BY_M9
`endif 

`ifdef i_axi_AXI_VV_S3_BY_M10
  `define AXI_VV_S3_BY_M10 `i_axi_AXI_VV_S3_BY_M10
`endif 

`ifdef i_axi_AXI_VV_S3_BY_M11
  `define AXI_VV_S3_BY_M11 `i_axi_AXI_VV_S3_BY_M11
`endif 

`ifdef i_axi_AXI_VV_S3_BY_M12
  `define AXI_VV_S3_BY_M12 `i_axi_AXI_VV_S3_BY_M12
`endif 

`ifdef i_axi_AXI_VV_S3_BY_M13
  `define AXI_VV_S3_BY_M13 `i_axi_AXI_VV_S3_BY_M13
`endif 

`ifdef i_axi_AXI_VV_S3_BY_M14
  `define AXI_VV_S3_BY_M14 `i_axi_AXI_VV_S3_BY_M14
`endif 

`ifdef i_axi_AXI_VV_S3_BY_M15
  `define AXI_VV_S3_BY_M15 `i_axi_AXI_VV_S3_BY_M15
`endif 

`ifdef i_axi_AXI_VV_S3_BY_M16
  `define AXI_VV_S3_BY_M16 `i_axi_AXI_VV_S3_BY_M16
`endif 

`ifdef i_axi_AXI_VV_S4_BY_M1
  `define AXI_VV_S4_BY_M1 `i_axi_AXI_VV_S4_BY_M1
`endif 

`ifdef i_axi_AXI_VV_S4_BY_M2
  `define AXI_VV_S4_BY_M2 `i_axi_AXI_VV_S4_BY_M2
`endif 

`ifdef i_axi_AXI_VV_S4_BY_M3
  `define AXI_VV_S4_BY_M3 `i_axi_AXI_VV_S4_BY_M3
`endif 

`ifdef i_axi_AXI_VV_S4_BY_M4
  `define AXI_VV_S4_BY_M4 `i_axi_AXI_VV_S4_BY_M4
`endif 

`ifdef i_axi_AXI_VV_S4_BY_M5
  `define AXI_VV_S4_BY_M5 `i_axi_AXI_VV_S4_BY_M5
`endif 

`ifdef i_axi_AXI_VV_S4_BY_M6
  `define AXI_VV_S4_BY_M6 `i_axi_AXI_VV_S4_BY_M6
`endif 

`ifdef i_axi_AXI_VV_S4_BY_M7
  `define AXI_VV_S4_BY_M7 `i_axi_AXI_VV_S4_BY_M7
`endif 

`ifdef i_axi_AXI_VV_S4_BY_M8
  `define AXI_VV_S4_BY_M8 `i_axi_AXI_VV_S4_BY_M8
`endif 

`ifdef i_axi_AXI_VV_S4_BY_M9
  `define AXI_VV_S4_BY_M9 `i_axi_AXI_VV_S4_BY_M9
`endif 

`ifdef i_axi_AXI_VV_S4_BY_M10
  `define AXI_VV_S4_BY_M10 `i_axi_AXI_VV_S4_BY_M10
`endif 

`ifdef i_axi_AXI_VV_S4_BY_M11
  `define AXI_VV_S4_BY_M11 `i_axi_AXI_VV_S4_BY_M11
`endif 

`ifdef i_axi_AXI_VV_S4_BY_M12
  `define AXI_VV_S4_BY_M12 `i_axi_AXI_VV_S4_BY_M12
`endif 

`ifdef i_axi_AXI_VV_S4_BY_M13
  `define AXI_VV_S4_BY_M13 `i_axi_AXI_VV_S4_BY_M13
`endif 

`ifdef i_axi_AXI_VV_S4_BY_M14
  `define AXI_VV_S4_BY_M14 `i_axi_AXI_VV_S4_BY_M14
`endif 

`ifdef i_axi_AXI_VV_S4_BY_M15
  `define AXI_VV_S4_BY_M15 `i_axi_AXI_VV_S4_BY_M15
`endif 

`ifdef i_axi_AXI_VV_S4_BY_M16
  `define AXI_VV_S4_BY_M16 `i_axi_AXI_VV_S4_BY_M16
`endif 

`ifdef i_axi_AXI_VV_S5_BY_M1
  `define AXI_VV_S5_BY_M1 `i_axi_AXI_VV_S5_BY_M1
`endif 

`ifdef i_axi_AXI_VV_S5_BY_M2
  `define AXI_VV_S5_BY_M2 `i_axi_AXI_VV_S5_BY_M2
`endif 

`ifdef i_axi_AXI_VV_S5_BY_M3
  `define AXI_VV_S5_BY_M3 `i_axi_AXI_VV_S5_BY_M3
`endif 

`ifdef i_axi_AXI_VV_S5_BY_M4
  `define AXI_VV_S5_BY_M4 `i_axi_AXI_VV_S5_BY_M4
`endif 

`ifdef i_axi_AXI_VV_S5_BY_M5
  `define AXI_VV_S5_BY_M5 `i_axi_AXI_VV_S5_BY_M5
`endif 

`ifdef i_axi_AXI_VV_S5_BY_M6
  `define AXI_VV_S5_BY_M6 `i_axi_AXI_VV_S5_BY_M6
`endif 

`ifdef i_axi_AXI_VV_S5_BY_M7
  `define AXI_VV_S5_BY_M7 `i_axi_AXI_VV_S5_BY_M7
`endif 

`ifdef i_axi_AXI_VV_S5_BY_M8
  `define AXI_VV_S5_BY_M8 `i_axi_AXI_VV_S5_BY_M8
`endif 

`ifdef i_axi_AXI_VV_S5_BY_M9
  `define AXI_VV_S5_BY_M9 `i_axi_AXI_VV_S5_BY_M9
`endif 

`ifdef i_axi_AXI_VV_S5_BY_M10
  `define AXI_VV_S5_BY_M10 `i_axi_AXI_VV_S5_BY_M10
`endif 

`ifdef i_axi_AXI_VV_S5_BY_M11
  `define AXI_VV_S5_BY_M11 `i_axi_AXI_VV_S5_BY_M11
`endif 

`ifdef i_axi_AXI_VV_S5_BY_M12
  `define AXI_VV_S5_BY_M12 `i_axi_AXI_VV_S5_BY_M12
`endif 

`ifdef i_axi_AXI_VV_S5_BY_M13
  `define AXI_VV_S5_BY_M13 `i_axi_AXI_VV_S5_BY_M13
`endif 

`ifdef i_axi_AXI_VV_S5_BY_M14
  `define AXI_VV_S5_BY_M14 `i_axi_AXI_VV_S5_BY_M14
`endif 

`ifdef i_axi_AXI_VV_S5_BY_M15
  `define AXI_VV_S5_BY_M15 `i_axi_AXI_VV_S5_BY_M15
`endif 

`ifdef i_axi_AXI_VV_S5_BY_M16
  `define AXI_VV_S5_BY_M16 `i_axi_AXI_VV_S5_BY_M16
`endif 

`ifdef i_axi_AXI_VV_S6_BY_M1
  `define AXI_VV_S6_BY_M1 `i_axi_AXI_VV_S6_BY_M1
`endif 

`ifdef i_axi_AXI_VV_S6_BY_M2
  `define AXI_VV_S6_BY_M2 `i_axi_AXI_VV_S6_BY_M2
`endif 

`ifdef i_axi_AXI_VV_S6_BY_M3
  `define AXI_VV_S6_BY_M3 `i_axi_AXI_VV_S6_BY_M3
`endif 

`ifdef i_axi_AXI_VV_S6_BY_M4
  `define AXI_VV_S6_BY_M4 `i_axi_AXI_VV_S6_BY_M4
`endif 

`ifdef i_axi_AXI_VV_S6_BY_M5
  `define AXI_VV_S6_BY_M5 `i_axi_AXI_VV_S6_BY_M5
`endif 

`ifdef i_axi_AXI_VV_S6_BY_M6
  `define AXI_VV_S6_BY_M6 `i_axi_AXI_VV_S6_BY_M6
`endif 

`ifdef i_axi_AXI_VV_S6_BY_M7
  `define AXI_VV_S6_BY_M7 `i_axi_AXI_VV_S6_BY_M7
`endif 

`ifdef i_axi_AXI_VV_S6_BY_M8
  `define AXI_VV_S6_BY_M8 `i_axi_AXI_VV_S6_BY_M8
`endif 

`ifdef i_axi_AXI_VV_S6_BY_M9
  `define AXI_VV_S6_BY_M9 `i_axi_AXI_VV_S6_BY_M9
`endif 

`ifdef i_axi_AXI_VV_S6_BY_M10
  `define AXI_VV_S6_BY_M10 `i_axi_AXI_VV_S6_BY_M10
`endif 

`ifdef i_axi_AXI_VV_S6_BY_M11
  `define AXI_VV_S6_BY_M11 `i_axi_AXI_VV_S6_BY_M11
`endif 

`ifdef i_axi_AXI_VV_S6_BY_M12
  `define AXI_VV_S6_BY_M12 `i_axi_AXI_VV_S6_BY_M12
`endif 

`ifdef i_axi_AXI_VV_S6_BY_M13
  `define AXI_VV_S6_BY_M13 `i_axi_AXI_VV_S6_BY_M13
`endif 

`ifdef i_axi_AXI_VV_S6_BY_M14
  `define AXI_VV_S6_BY_M14 `i_axi_AXI_VV_S6_BY_M14
`endif 

`ifdef i_axi_AXI_VV_S6_BY_M15
  `define AXI_VV_S6_BY_M15 `i_axi_AXI_VV_S6_BY_M15
`endif 

`ifdef i_axi_AXI_VV_S6_BY_M16
  `define AXI_VV_S6_BY_M16 `i_axi_AXI_VV_S6_BY_M16
`endif 

`ifdef i_axi_AXI_VV_S7_BY_M1
  `define AXI_VV_S7_BY_M1 `i_axi_AXI_VV_S7_BY_M1
`endif 

`ifdef i_axi_AXI_VV_S7_BY_M2
  `define AXI_VV_S7_BY_M2 `i_axi_AXI_VV_S7_BY_M2
`endif 

`ifdef i_axi_AXI_VV_S7_BY_M3
  `define AXI_VV_S7_BY_M3 `i_axi_AXI_VV_S7_BY_M3
`endif 

`ifdef i_axi_AXI_VV_S7_BY_M4
  `define AXI_VV_S7_BY_M4 `i_axi_AXI_VV_S7_BY_M4
`endif 

`ifdef i_axi_AXI_VV_S7_BY_M5
  `define AXI_VV_S7_BY_M5 `i_axi_AXI_VV_S7_BY_M5
`endif 

`ifdef i_axi_AXI_VV_S7_BY_M6
  `define AXI_VV_S7_BY_M6 `i_axi_AXI_VV_S7_BY_M6
`endif 

`ifdef i_axi_AXI_VV_S7_BY_M7
  `define AXI_VV_S7_BY_M7 `i_axi_AXI_VV_S7_BY_M7
`endif 

`ifdef i_axi_AXI_VV_S7_BY_M8
  `define AXI_VV_S7_BY_M8 `i_axi_AXI_VV_S7_BY_M8
`endif 

`ifdef i_axi_AXI_VV_S7_BY_M9
  `define AXI_VV_S7_BY_M9 `i_axi_AXI_VV_S7_BY_M9
`endif 

`ifdef i_axi_AXI_VV_S7_BY_M10
  `define AXI_VV_S7_BY_M10 `i_axi_AXI_VV_S7_BY_M10
`endif 

`ifdef i_axi_AXI_VV_S7_BY_M11
  `define AXI_VV_S7_BY_M11 `i_axi_AXI_VV_S7_BY_M11
`endif 

`ifdef i_axi_AXI_VV_S7_BY_M12
  `define AXI_VV_S7_BY_M12 `i_axi_AXI_VV_S7_BY_M12
`endif 

`ifdef i_axi_AXI_VV_S7_BY_M13
  `define AXI_VV_S7_BY_M13 `i_axi_AXI_VV_S7_BY_M13
`endif 

`ifdef i_axi_AXI_VV_S7_BY_M14
  `define AXI_VV_S7_BY_M14 `i_axi_AXI_VV_S7_BY_M14
`endif 

`ifdef i_axi_AXI_VV_S7_BY_M15
  `define AXI_VV_S7_BY_M15 `i_axi_AXI_VV_S7_BY_M15
`endif 

`ifdef i_axi_AXI_VV_S7_BY_M16
  `define AXI_VV_S7_BY_M16 `i_axi_AXI_VV_S7_BY_M16
`endif 

`ifdef i_axi_AXI_VV_S8_BY_M1
  `define AXI_VV_S8_BY_M1 `i_axi_AXI_VV_S8_BY_M1
`endif 

`ifdef i_axi_AXI_VV_S8_BY_M2
  `define AXI_VV_S8_BY_M2 `i_axi_AXI_VV_S8_BY_M2
`endif 

`ifdef i_axi_AXI_VV_S8_BY_M3
  `define AXI_VV_S8_BY_M3 `i_axi_AXI_VV_S8_BY_M3
`endif 

`ifdef i_axi_AXI_VV_S8_BY_M4
  `define AXI_VV_S8_BY_M4 `i_axi_AXI_VV_S8_BY_M4
`endif 

`ifdef i_axi_AXI_VV_S8_BY_M5
  `define AXI_VV_S8_BY_M5 `i_axi_AXI_VV_S8_BY_M5
`endif 

`ifdef i_axi_AXI_VV_S8_BY_M6
  `define AXI_VV_S8_BY_M6 `i_axi_AXI_VV_S8_BY_M6
`endif 

`ifdef i_axi_AXI_VV_S8_BY_M7
  `define AXI_VV_S8_BY_M7 `i_axi_AXI_VV_S8_BY_M7
`endif 

`ifdef i_axi_AXI_VV_S8_BY_M8
  `define AXI_VV_S8_BY_M8 `i_axi_AXI_VV_S8_BY_M8
`endif 

`ifdef i_axi_AXI_VV_S8_BY_M9
  `define AXI_VV_S8_BY_M9 `i_axi_AXI_VV_S8_BY_M9
`endif 

`ifdef i_axi_AXI_VV_S8_BY_M10
  `define AXI_VV_S8_BY_M10 `i_axi_AXI_VV_S8_BY_M10
`endif 

`ifdef i_axi_AXI_VV_S8_BY_M11
  `define AXI_VV_S8_BY_M11 `i_axi_AXI_VV_S8_BY_M11
`endif 

`ifdef i_axi_AXI_VV_S8_BY_M12
  `define AXI_VV_S8_BY_M12 `i_axi_AXI_VV_S8_BY_M12
`endif 

`ifdef i_axi_AXI_VV_S8_BY_M13
  `define AXI_VV_S8_BY_M13 `i_axi_AXI_VV_S8_BY_M13
`endif 

`ifdef i_axi_AXI_VV_S8_BY_M14
  `define AXI_VV_S8_BY_M14 `i_axi_AXI_VV_S8_BY_M14
`endif 

`ifdef i_axi_AXI_VV_S8_BY_M15
  `define AXI_VV_S8_BY_M15 `i_axi_AXI_VV_S8_BY_M15
`endif 

`ifdef i_axi_AXI_VV_S8_BY_M16
  `define AXI_VV_S8_BY_M16 `i_axi_AXI_VV_S8_BY_M16
`endif 

`ifdef i_axi_AXI_VV_S9_BY_M1
  `define AXI_VV_S9_BY_M1 `i_axi_AXI_VV_S9_BY_M1
`endif 

`ifdef i_axi_AXI_VV_S9_BY_M2
  `define AXI_VV_S9_BY_M2 `i_axi_AXI_VV_S9_BY_M2
`endif 

`ifdef i_axi_AXI_VV_S9_BY_M3
  `define AXI_VV_S9_BY_M3 `i_axi_AXI_VV_S9_BY_M3
`endif 

`ifdef i_axi_AXI_VV_S9_BY_M4
  `define AXI_VV_S9_BY_M4 `i_axi_AXI_VV_S9_BY_M4
`endif 

`ifdef i_axi_AXI_VV_S9_BY_M5
  `define AXI_VV_S9_BY_M5 `i_axi_AXI_VV_S9_BY_M5
`endif 

`ifdef i_axi_AXI_VV_S9_BY_M6
  `define AXI_VV_S9_BY_M6 `i_axi_AXI_VV_S9_BY_M6
`endif 

`ifdef i_axi_AXI_VV_S9_BY_M7
  `define AXI_VV_S9_BY_M7 `i_axi_AXI_VV_S9_BY_M7
`endif 

`ifdef i_axi_AXI_VV_S9_BY_M8
  `define AXI_VV_S9_BY_M8 `i_axi_AXI_VV_S9_BY_M8
`endif 

`ifdef i_axi_AXI_VV_S9_BY_M9
  `define AXI_VV_S9_BY_M9 `i_axi_AXI_VV_S9_BY_M9
`endif 

`ifdef i_axi_AXI_VV_S9_BY_M10
  `define AXI_VV_S9_BY_M10 `i_axi_AXI_VV_S9_BY_M10
`endif 

`ifdef i_axi_AXI_VV_S9_BY_M11
  `define AXI_VV_S9_BY_M11 `i_axi_AXI_VV_S9_BY_M11
`endif 

`ifdef i_axi_AXI_VV_S9_BY_M12
  `define AXI_VV_S9_BY_M12 `i_axi_AXI_VV_S9_BY_M12
`endif 

`ifdef i_axi_AXI_VV_S9_BY_M13
  `define AXI_VV_S9_BY_M13 `i_axi_AXI_VV_S9_BY_M13
`endif 

`ifdef i_axi_AXI_VV_S9_BY_M14
  `define AXI_VV_S9_BY_M14 `i_axi_AXI_VV_S9_BY_M14
`endif 

`ifdef i_axi_AXI_VV_S9_BY_M15
  `define AXI_VV_S9_BY_M15 `i_axi_AXI_VV_S9_BY_M15
`endif 

`ifdef i_axi_AXI_VV_S9_BY_M16
  `define AXI_VV_S9_BY_M16 `i_axi_AXI_VV_S9_BY_M16
`endif 

`ifdef i_axi_AXI_VV_S10_BY_M1
  `define AXI_VV_S10_BY_M1 `i_axi_AXI_VV_S10_BY_M1
`endif 

`ifdef i_axi_AXI_VV_S10_BY_M2
  `define AXI_VV_S10_BY_M2 `i_axi_AXI_VV_S10_BY_M2
`endif 

`ifdef i_axi_AXI_VV_S10_BY_M3
  `define AXI_VV_S10_BY_M3 `i_axi_AXI_VV_S10_BY_M3
`endif 

`ifdef i_axi_AXI_VV_S10_BY_M4
  `define AXI_VV_S10_BY_M4 `i_axi_AXI_VV_S10_BY_M4
`endif 

`ifdef i_axi_AXI_VV_S10_BY_M5
  `define AXI_VV_S10_BY_M5 `i_axi_AXI_VV_S10_BY_M5
`endif 

`ifdef i_axi_AXI_VV_S10_BY_M6
  `define AXI_VV_S10_BY_M6 `i_axi_AXI_VV_S10_BY_M6
`endif 

`ifdef i_axi_AXI_VV_S10_BY_M7
  `define AXI_VV_S10_BY_M7 `i_axi_AXI_VV_S10_BY_M7
`endif 

`ifdef i_axi_AXI_VV_S10_BY_M8
  `define AXI_VV_S10_BY_M8 `i_axi_AXI_VV_S10_BY_M8
`endif 

`ifdef i_axi_AXI_VV_S10_BY_M9
  `define AXI_VV_S10_BY_M9 `i_axi_AXI_VV_S10_BY_M9
`endif 

`ifdef i_axi_AXI_VV_S10_BY_M10
  `define AXI_VV_S10_BY_M10 `i_axi_AXI_VV_S10_BY_M10
`endif 

`ifdef i_axi_AXI_VV_S10_BY_M11
  `define AXI_VV_S10_BY_M11 `i_axi_AXI_VV_S10_BY_M11
`endif 

`ifdef i_axi_AXI_VV_S10_BY_M12
  `define AXI_VV_S10_BY_M12 `i_axi_AXI_VV_S10_BY_M12
`endif 

`ifdef i_axi_AXI_VV_S10_BY_M13
  `define AXI_VV_S10_BY_M13 `i_axi_AXI_VV_S10_BY_M13
`endif 

`ifdef i_axi_AXI_VV_S10_BY_M14
  `define AXI_VV_S10_BY_M14 `i_axi_AXI_VV_S10_BY_M14
`endif 

`ifdef i_axi_AXI_VV_S10_BY_M15
  `define AXI_VV_S10_BY_M15 `i_axi_AXI_VV_S10_BY_M15
`endif 

`ifdef i_axi_AXI_VV_S10_BY_M16
  `define AXI_VV_S10_BY_M16 `i_axi_AXI_VV_S10_BY_M16
`endif 

`ifdef i_axi_AXI_VV_S11_BY_M1
  `define AXI_VV_S11_BY_M1 `i_axi_AXI_VV_S11_BY_M1
`endif 

`ifdef i_axi_AXI_VV_S11_BY_M2
  `define AXI_VV_S11_BY_M2 `i_axi_AXI_VV_S11_BY_M2
`endif 

`ifdef i_axi_AXI_VV_S11_BY_M3
  `define AXI_VV_S11_BY_M3 `i_axi_AXI_VV_S11_BY_M3
`endif 

`ifdef i_axi_AXI_VV_S11_BY_M4
  `define AXI_VV_S11_BY_M4 `i_axi_AXI_VV_S11_BY_M4
`endif 

`ifdef i_axi_AXI_VV_S11_BY_M5
  `define AXI_VV_S11_BY_M5 `i_axi_AXI_VV_S11_BY_M5
`endif 

`ifdef i_axi_AXI_VV_S11_BY_M6
  `define AXI_VV_S11_BY_M6 `i_axi_AXI_VV_S11_BY_M6
`endif 

`ifdef i_axi_AXI_VV_S11_BY_M7
  `define AXI_VV_S11_BY_M7 `i_axi_AXI_VV_S11_BY_M7
`endif 

`ifdef i_axi_AXI_VV_S11_BY_M8
  `define AXI_VV_S11_BY_M8 `i_axi_AXI_VV_S11_BY_M8
`endif 

`ifdef i_axi_AXI_VV_S11_BY_M9
  `define AXI_VV_S11_BY_M9 `i_axi_AXI_VV_S11_BY_M9
`endif 

`ifdef i_axi_AXI_VV_S11_BY_M10
  `define AXI_VV_S11_BY_M10 `i_axi_AXI_VV_S11_BY_M10
`endif 

`ifdef i_axi_AXI_VV_S11_BY_M11
  `define AXI_VV_S11_BY_M11 `i_axi_AXI_VV_S11_BY_M11
`endif 

`ifdef i_axi_AXI_VV_S11_BY_M12
  `define AXI_VV_S11_BY_M12 `i_axi_AXI_VV_S11_BY_M12
`endif 

`ifdef i_axi_AXI_VV_S11_BY_M13
  `define AXI_VV_S11_BY_M13 `i_axi_AXI_VV_S11_BY_M13
`endif 

`ifdef i_axi_AXI_VV_S11_BY_M14
  `define AXI_VV_S11_BY_M14 `i_axi_AXI_VV_S11_BY_M14
`endif 

`ifdef i_axi_AXI_VV_S11_BY_M15
  `define AXI_VV_S11_BY_M15 `i_axi_AXI_VV_S11_BY_M15
`endif 

`ifdef i_axi_AXI_VV_S11_BY_M16
  `define AXI_VV_S11_BY_M16 `i_axi_AXI_VV_S11_BY_M16
`endif 

`ifdef i_axi_AXI_VV_S12_BY_M1
  `define AXI_VV_S12_BY_M1 `i_axi_AXI_VV_S12_BY_M1
`endif 

`ifdef i_axi_AXI_VV_S12_BY_M2
  `define AXI_VV_S12_BY_M2 `i_axi_AXI_VV_S12_BY_M2
`endif 

`ifdef i_axi_AXI_VV_S12_BY_M3
  `define AXI_VV_S12_BY_M3 `i_axi_AXI_VV_S12_BY_M3
`endif 

`ifdef i_axi_AXI_VV_S12_BY_M4
  `define AXI_VV_S12_BY_M4 `i_axi_AXI_VV_S12_BY_M4
`endif 

`ifdef i_axi_AXI_VV_S12_BY_M5
  `define AXI_VV_S12_BY_M5 `i_axi_AXI_VV_S12_BY_M5
`endif 

`ifdef i_axi_AXI_VV_S12_BY_M6
  `define AXI_VV_S12_BY_M6 `i_axi_AXI_VV_S12_BY_M6
`endif 

`ifdef i_axi_AXI_VV_S12_BY_M7
  `define AXI_VV_S12_BY_M7 `i_axi_AXI_VV_S12_BY_M7
`endif 

`ifdef i_axi_AXI_VV_S12_BY_M8
  `define AXI_VV_S12_BY_M8 `i_axi_AXI_VV_S12_BY_M8
`endif 

`ifdef i_axi_AXI_VV_S12_BY_M9
  `define AXI_VV_S12_BY_M9 `i_axi_AXI_VV_S12_BY_M9
`endif 

`ifdef i_axi_AXI_VV_S12_BY_M10
  `define AXI_VV_S12_BY_M10 `i_axi_AXI_VV_S12_BY_M10
`endif 

`ifdef i_axi_AXI_VV_S12_BY_M11
  `define AXI_VV_S12_BY_M11 `i_axi_AXI_VV_S12_BY_M11
`endif 

`ifdef i_axi_AXI_VV_S12_BY_M12
  `define AXI_VV_S12_BY_M12 `i_axi_AXI_VV_S12_BY_M12
`endif 

`ifdef i_axi_AXI_VV_S12_BY_M13
  `define AXI_VV_S12_BY_M13 `i_axi_AXI_VV_S12_BY_M13
`endif 

`ifdef i_axi_AXI_VV_S12_BY_M14
  `define AXI_VV_S12_BY_M14 `i_axi_AXI_VV_S12_BY_M14
`endif 

`ifdef i_axi_AXI_VV_S12_BY_M15
  `define AXI_VV_S12_BY_M15 `i_axi_AXI_VV_S12_BY_M15
`endif 

`ifdef i_axi_AXI_VV_S12_BY_M16
  `define AXI_VV_S12_BY_M16 `i_axi_AXI_VV_S12_BY_M16
`endif 

`ifdef i_axi_AXI_VV_S13_BY_M1
  `define AXI_VV_S13_BY_M1 `i_axi_AXI_VV_S13_BY_M1
`endif 

`ifdef i_axi_AXI_VV_S13_BY_M2
  `define AXI_VV_S13_BY_M2 `i_axi_AXI_VV_S13_BY_M2
`endif 

`ifdef i_axi_AXI_VV_S13_BY_M3
  `define AXI_VV_S13_BY_M3 `i_axi_AXI_VV_S13_BY_M3
`endif 

`ifdef i_axi_AXI_VV_S13_BY_M4
  `define AXI_VV_S13_BY_M4 `i_axi_AXI_VV_S13_BY_M4
`endif 

`ifdef i_axi_AXI_VV_S13_BY_M5
  `define AXI_VV_S13_BY_M5 `i_axi_AXI_VV_S13_BY_M5
`endif 

`ifdef i_axi_AXI_VV_S13_BY_M6
  `define AXI_VV_S13_BY_M6 `i_axi_AXI_VV_S13_BY_M6
`endif 

`ifdef i_axi_AXI_VV_S13_BY_M7
  `define AXI_VV_S13_BY_M7 `i_axi_AXI_VV_S13_BY_M7
`endif 

`ifdef i_axi_AXI_VV_S13_BY_M8
  `define AXI_VV_S13_BY_M8 `i_axi_AXI_VV_S13_BY_M8
`endif 

`ifdef i_axi_AXI_VV_S13_BY_M9
  `define AXI_VV_S13_BY_M9 `i_axi_AXI_VV_S13_BY_M9
`endif 

`ifdef i_axi_AXI_VV_S13_BY_M10
  `define AXI_VV_S13_BY_M10 `i_axi_AXI_VV_S13_BY_M10
`endif 

`ifdef i_axi_AXI_VV_S13_BY_M11
  `define AXI_VV_S13_BY_M11 `i_axi_AXI_VV_S13_BY_M11
`endif 

`ifdef i_axi_AXI_VV_S13_BY_M12
  `define AXI_VV_S13_BY_M12 `i_axi_AXI_VV_S13_BY_M12
`endif 

`ifdef i_axi_AXI_VV_S13_BY_M13
  `define AXI_VV_S13_BY_M13 `i_axi_AXI_VV_S13_BY_M13
`endif 

`ifdef i_axi_AXI_VV_S13_BY_M14
  `define AXI_VV_S13_BY_M14 `i_axi_AXI_VV_S13_BY_M14
`endif 

`ifdef i_axi_AXI_VV_S13_BY_M15
  `define AXI_VV_S13_BY_M15 `i_axi_AXI_VV_S13_BY_M15
`endif 

`ifdef i_axi_AXI_VV_S13_BY_M16
  `define AXI_VV_S13_BY_M16 `i_axi_AXI_VV_S13_BY_M16
`endif 

`ifdef i_axi_AXI_VV_S14_BY_M1
  `define AXI_VV_S14_BY_M1 `i_axi_AXI_VV_S14_BY_M1
`endif 

`ifdef i_axi_AXI_VV_S14_BY_M2
  `define AXI_VV_S14_BY_M2 `i_axi_AXI_VV_S14_BY_M2
`endif 

`ifdef i_axi_AXI_VV_S14_BY_M3
  `define AXI_VV_S14_BY_M3 `i_axi_AXI_VV_S14_BY_M3
`endif 

`ifdef i_axi_AXI_VV_S14_BY_M4
  `define AXI_VV_S14_BY_M4 `i_axi_AXI_VV_S14_BY_M4
`endif 

`ifdef i_axi_AXI_VV_S14_BY_M5
  `define AXI_VV_S14_BY_M5 `i_axi_AXI_VV_S14_BY_M5
`endif 

`ifdef i_axi_AXI_VV_S14_BY_M6
  `define AXI_VV_S14_BY_M6 `i_axi_AXI_VV_S14_BY_M6
`endif 

`ifdef i_axi_AXI_VV_S14_BY_M7
  `define AXI_VV_S14_BY_M7 `i_axi_AXI_VV_S14_BY_M7
`endif 

`ifdef i_axi_AXI_VV_S14_BY_M8
  `define AXI_VV_S14_BY_M8 `i_axi_AXI_VV_S14_BY_M8
`endif 

`ifdef i_axi_AXI_VV_S14_BY_M9
  `define AXI_VV_S14_BY_M9 `i_axi_AXI_VV_S14_BY_M9
`endif 

`ifdef i_axi_AXI_VV_S14_BY_M10
  `define AXI_VV_S14_BY_M10 `i_axi_AXI_VV_S14_BY_M10
`endif 

`ifdef i_axi_AXI_VV_S14_BY_M11
  `define AXI_VV_S14_BY_M11 `i_axi_AXI_VV_S14_BY_M11
`endif 

`ifdef i_axi_AXI_VV_S14_BY_M12
  `define AXI_VV_S14_BY_M12 `i_axi_AXI_VV_S14_BY_M12
`endif 

`ifdef i_axi_AXI_VV_S14_BY_M13
  `define AXI_VV_S14_BY_M13 `i_axi_AXI_VV_S14_BY_M13
`endif 

`ifdef i_axi_AXI_VV_S14_BY_M14
  `define AXI_VV_S14_BY_M14 `i_axi_AXI_VV_S14_BY_M14
`endif 

`ifdef i_axi_AXI_VV_S14_BY_M15
  `define AXI_VV_S14_BY_M15 `i_axi_AXI_VV_S14_BY_M15
`endif 

`ifdef i_axi_AXI_VV_S14_BY_M16
  `define AXI_VV_S14_BY_M16 `i_axi_AXI_VV_S14_BY_M16
`endif 

`ifdef i_axi_AXI_VV_S15_BY_M1
  `define AXI_VV_S15_BY_M1 `i_axi_AXI_VV_S15_BY_M1
`endif 

`ifdef i_axi_AXI_VV_S15_BY_M2
  `define AXI_VV_S15_BY_M2 `i_axi_AXI_VV_S15_BY_M2
`endif 

`ifdef i_axi_AXI_VV_S15_BY_M3
  `define AXI_VV_S15_BY_M3 `i_axi_AXI_VV_S15_BY_M3
`endif 

`ifdef i_axi_AXI_VV_S15_BY_M4
  `define AXI_VV_S15_BY_M4 `i_axi_AXI_VV_S15_BY_M4
`endif 

`ifdef i_axi_AXI_VV_S15_BY_M5
  `define AXI_VV_S15_BY_M5 `i_axi_AXI_VV_S15_BY_M5
`endif 

`ifdef i_axi_AXI_VV_S15_BY_M6
  `define AXI_VV_S15_BY_M6 `i_axi_AXI_VV_S15_BY_M6
`endif 

`ifdef i_axi_AXI_VV_S15_BY_M7
  `define AXI_VV_S15_BY_M7 `i_axi_AXI_VV_S15_BY_M7
`endif 

`ifdef i_axi_AXI_VV_S15_BY_M8
  `define AXI_VV_S15_BY_M8 `i_axi_AXI_VV_S15_BY_M8
`endif 

`ifdef i_axi_AXI_VV_S15_BY_M9
  `define AXI_VV_S15_BY_M9 `i_axi_AXI_VV_S15_BY_M9
`endif 

`ifdef i_axi_AXI_VV_S15_BY_M10
  `define AXI_VV_S15_BY_M10 `i_axi_AXI_VV_S15_BY_M10
`endif 

`ifdef i_axi_AXI_VV_S15_BY_M11
  `define AXI_VV_S15_BY_M11 `i_axi_AXI_VV_S15_BY_M11
`endif 

`ifdef i_axi_AXI_VV_S15_BY_M12
  `define AXI_VV_S15_BY_M12 `i_axi_AXI_VV_S15_BY_M12
`endif 

`ifdef i_axi_AXI_VV_S15_BY_M13
  `define AXI_VV_S15_BY_M13 `i_axi_AXI_VV_S15_BY_M13
`endif 

`ifdef i_axi_AXI_VV_S15_BY_M14
  `define AXI_VV_S15_BY_M14 `i_axi_AXI_VV_S15_BY_M14
`endif 

`ifdef i_axi_AXI_VV_S15_BY_M15
  `define AXI_VV_S15_BY_M15 `i_axi_AXI_VV_S15_BY_M15
`endif 

`ifdef i_axi_AXI_VV_S15_BY_M16
  `define AXI_VV_S15_BY_M16 `i_axi_AXI_VV_S15_BY_M16
`endif 

`ifdef i_axi_AXI_VV_S16_BY_M1
  `define AXI_VV_S16_BY_M1 `i_axi_AXI_VV_S16_BY_M1
`endif 

`ifdef i_axi_AXI_VV_S16_BY_M2
  `define AXI_VV_S16_BY_M2 `i_axi_AXI_VV_S16_BY_M2
`endif 

`ifdef i_axi_AXI_VV_S16_BY_M3
  `define AXI_VV_S16_BY_M3 `i_axi_AXI_VV_S16_BY_M3
`endif 

`ifdef i_axi_AXI_VV_S16_BY_M4
  `define AXI_VV_S16_BY_M4 `i_axi_AXI_VV_S16_BY_M4
`endif 

`ifdef i_axi_AXI_VV_S16_BY_M5
  `define AXI_VV_S16_BY_M5 `i_axi_AXI_VV_S16_BY_M5
`endif 

`ifdef i_axi_AXI_VV_S16_BY_M6
  `define AXI_VV_S16_BY_M6 `i_axi_AXI_VV_S16_BY_M6
`endif 

`ifdef i_axi_AXI_VV_S16_BY_M7
  `define AXI_VV_S16_BY_M7 `i_axi_AXI_VV_S16_BY_M7
`endif 

`ifdef i_axi_AXI_VV_S16_BY_M8
  `define AXI_VV_S16_BY_M8 `i_axi_AXI_VV_S16_BY_M8
`endif 

`ifdef i_axi_AXI_VV_S16_BY_M9
  `define AXI_VV_S16_BY_M9 `i_axi_AXI_VV_S16_BY_M9
`endif 

`ifdef i_axi_AXI_VV_S16_BY_M10
  `define AXI_VV_S16_BY_M10 `i_axi_AXI_VV_S16_BY_M10
`endif 

`ifdef i_axi_AXI_VV_S16_BY_M11
  `define AXI_VV_S16_BY_M11 `i_axi_AXI_VV_S16_BY_M11
`endif 

`ifdef i_axi_AXI_VV_S16_BY_M12
  `define AXI_VV_S16_BY_M12 `i_axi_AXI_VV_S16_BY_M12
`endif 

`ifdef i_axi_AXI_VV_S16_BY_M13
  `define AXI_VV_S16_BY_M13 `i_axi_AXI_VV_S16_BY_M13
`endif 

`ifdef i_axi_AXI_VV_S16_BY_M14
  `define AXI_VV_S16_BY_M14 `i_axi_AXI_VV_S16_BY_M14
`endif 

`ifdef i_axi_AXI_VV_S16_BY_M15
  `define AXI_VV_S16_BY_M15 `i_axi_AXI_VV_S16_BY_M15
`endif 

`ifdef i_axi_AXI_VV_S16_BY_M16
  `define AXI_VV_S16_BY_M16 `i_axi_AXI_VV_S16_BY_M16
`endif 

`ifdef i_axi_AXI_NMV_S1
  `define AXI_NMV_S1 `i_axi_AXI_NMV_S1
`endif 

`ifdef i_axi_AXI_LOG2_NMV_S1
  `define AXI_LOG2_NMV_S1 `i_axi_AXI_LOG2_NMV_S1
`endif 

`ifdef i_axi_AXI_LOG2_NMP1V_S1
  `define AXI_LOG2_NMP1V_S1 `i_axi_AXI_LOG2_NMP1V_S1
`endif 

`ifdef i_axi_AXI_NMV_S2
  `define AXI_NMV_S2 `i_axi_AXI_NMV_S2
`endif 

`ifdef i_axi_AXI_LOG2_NMV_S2
  `define AXI_LOG2_NMV_S2 `i_axi_AXI_LOG2_NMV_S2
`endif 

`ifdef i_axi_AXI_LOG2_NMP1V_S2
  `define AXI_LOG2_NMP1V_S2 `i_axi_AXI_LOG2_NMP1V_S2
`endif 

`ifdef i_axi_AXI_NMV_S3
  `define AXI_NMV_S3 `i_axi_AXI_NMV_S3
`endif 

`ifdef i_axi_AXI_LOG2_NMV_S3
  `define AXI_LOG2_NMV_S3 `i_axi_AXI_LOG2_NMV_S3
`endif 

`ifdef i_axi_AXI_LOG2_NMP1V_S3
  `define AXI_LOG2_NMP1V_S3 `i_axi_AXI_LOG2_NMP1V_S3
`endif 

`ifdef i_axi_AXI_NMV_S4
  `define AXI_NMV_S4 `i_axi_AXI_NMV_S4
`endif 

`ifdef i_axi_AXI_LOG2_NMV_S4
  `define AXI_LOG2_NMV_S4 `i_axi_AXI_LOG2_NMV_S4
`endif 

`ifdef i_axi_AXI_LOG2_NMP1V_S4
  `define AXI_LOG2_NMP1V_S4 `i_axi_AXI_LOG2_NMP1V_S4
`endif 

`ifdef i_axi_AXI_NMV_S5
  `define AXI_NMV_S5 `i_axi_AXI_NMV_S5
`endif 

`ifdef i_axi_AXI_LOG2_NMV_S5
  `define AXI_LOG2_NMV_S5 `i_axi_AXI_LOG2_NMV_S5
`endif 

`ifdef i_axi_AXI_LOG2_NMP1V_S5
  `define AXI_LOG2_NMP1V_S5 `i_axi_AXI_LOG2_NMP1V_S5
`endif 

`ifdef i_axi_AXI_NMV_S6
  `define AXI_NMV_S6 `i_axi_AXI_NMV_S6
`endif 

`ifdef i_axi_AXI_LOG2_NMV_S6
  `define AXI_LOG2_NMV_S6 `i_axi_AXI_LOG2_NMV_S6
`endif 

`ifdef i_axi_AXI_LOG2_NMP1V_S6
  `define AXI_LOG2_NMP1V_S6 `i_axi_AXI_LOG2_NMP1V_S6
`endif 

`ifdef i_axi_AXI_NMV_S7
  `define AXI_NMV_S7 `i_axi_AXI_NMV_S7
`endif 

`ifdef i_axi_AXI_LOG2_NMV_S7
  `define AXI_LOG2_NMV_S7 `i_axi_AXI_LOG2_NMV_S7
`endif 

`ifdef i_axi_AXI_LOG2_NMP1V_S7
  `define AXI_LOG2_NMP1V_S7 `i_axi_AXI_LOG2_NMP1V_S7
`endif 

`ifdef i_axi_AXI_NMV_S8
  `define AXI_NMV_S8 `i_axi_AXI_NMV_S8
`endif 

`ifdef i_axi_AXI_LOG2_NMV_S8
  `define AXI_LOG2_NMV_S8 `i_axi_AXI_LOG2_NMV_S8
`endif 

`ifdef i_axi_AXI_LOG2_NMP1V_S8
  `define AXI_LOG2_NMP1V_S8 `i_axi_AXI_LOG2_NMP1V_S8
`endif 

`ifdef i_axi_AXI_NMV_S9
  `define AXI_NMV_S9 `i_axi_AXI_NMV_S9
`endif 

`ifdef i_axi_AXI_LOG2_NMV_S9
  `define AXI_LOG2_NMV_S9 `i_axi_AXI_LOG2_NMV_S9
`endif 

`ifdef i_axi_AXI_LOG2_NMP1V_S9
  `define AXI_LOG2_NMP1V_S9 `i_axi_AXI_LOG2_NMP1V_S9
`endif 

`ifdef i_axi_AXI_NMV_S10
  `define AXI_NMV_S10 `i_axi_AXI_NMV_S10
`endif 

`ifdef i_axi_AXI_LOG2_NMV_S10
  `define AXI_LOG2_NMV_S10 `i_axi_AXI_LOG2_NMV_S10
`endif 

`ifdef i_axi_AXI_LOG2_NMP1V_S10
  `define AXI_LOG2_NMP1V_S10 `i_axi_AXI_LOG2_NMP1V_S10
`endif 

`ifdef i_axi_AXI_NMV_S11
  `define AXI_NMV_S11 `i_axi_AXI_NMV_S11
`endif 

`ifdef i_axi_AXI_LOG2_NMV_S11
  `define AXI_LOG2_NMV_S11 `i_axi_AXI_LOG2_NMV_S11
`endif 

`ifdef i_axi_AXI_LOG2_NMP1V_S11
  `define AXI_LOG2_NMP1V_S11 `i_axi_AXI_LOG2_NMP1V_S11
`endif 

`ifdef i_axi_AXI_NMV_S12
  `define AXI_NMV_S12 `i_axi_AXI_NMV_S12
`endif 

`ifdef i_axi_AXI_LOG2_NMV_S12
  `define AXI_LOG2_NMV_S12 `i_axi_AXI_LOG2_NMV_S12
`endif 

`ifdef i_axi_AXI_LOG2_NMP1V_S12
  `define AXI_LOG2_NMP1V_S12 `i_axi_AXI_LOG2_NMP1V_S12
`endif 

`ifdef i_axi_AXI_NMV_S13
  `define AXI_NMV_S13 `i_axi_AXI_NMV_S13
`endif 

`ifdef i_axi_AXI_LOG2_NMV_S13
  `define AXI_LOG2_NMV_S13 `i_axi_AXI_LOG2_NMV_S13
`endif 

`ifdef i_axi_AXI_LOG2_NMP1V_S13
  `define AXI_LOG2_NMP1V_S13 `i_axi_AXI_LOG2_NMP1V_S13
`endif 

`ifdef i_axi_AXI_NMV_S14
  `define AXI_NMV_S14 `i_axi_AXI_NMV_S14
`endif 

`ifdef i_axi_AXI_LOG2_NMV_S14
  `define AXI_LOG2_NMV_S14 `i_axi_AXI_LOG2_NMV_S14
`endif 

`ifdef i_axi_AXI_LOG2_NMP1V_S14
  `define AXI_LOG2_NMP1V_S14 `i_axi_AXI_LOG2_NMP1V_S14
`endif 

`ifdef i_axi_AXI_NMV_S15
  `define AXI_NMV_S15 `i_axi_AXI_NMV_S15
`endif 

`ifdef i_axi_AXI_LOG2_NMV_S15
  `define AXI_LOG2_NMV_S15 `i_axi_AXI_LOG2_NMV_S15
`endif 

`ifdef i_axi_AXI_LOG2_NMP1V_S15
  `define AXI_LOG2_NMP1V_S15 `i_axi_AXI_LOG2_NMP1V_S15
`endif 

`ifdef i_axi_AXI_NMV_S16
  `define AXI_NMV_S16 `i_axi_AXI_NMV_S16
`endif 

`ifdef i_axi_AXI_LOG2_NMV_S16
  `define AXI_LOG2_NMV_S16 `i_axi_AXI_LOG2_NMV_S16
`endif 

`ifdef i_axi_AXI_LOG2_NMP1V_S16
  `define AXI_LOG2_NMP1V_S16 `i_axi_AXI_LOG2_NMP1V_S16
`endif 

`ifdef i_axi_AXI_NSV_M1
  `define AXI_NSV_M1 `i_axi_AXI_NSV_M1
`endif 

`ifdef i_axi_AXI_LOG2_NSV_M1
  `define AXI_LOG2_NSV_M1 `i_axi_AXI_LOG2_NSV_M1
`endif 

`ifdef i_axi_AXI_NSV_M2
  `define AXI_NSV_M2 `i_axi_AXI_NSV_M2
`endif 

`ifdef i_axi_AXI_LOG2_NSV_M2
  `define AXI_LOG2_NSV_M2 `i_axi_AXI_LOG2_NSV_M2
`endif 

`ifdef i_axi_AXI_NSV_M3
  `define AXI_NSV_M3 `i_axi_AXI_NSV_M3
`endif 

`ifdef i_axi_AXI_LOG2_NSV_M3
  `define AXI_LOG2_NSV_M3 `i_axi_AXI_LOG2_NSV_M3
`endif 

`ifdef i_axi_AXI_NSV_M4
  `define AXI_NSV_M4 `i_axi_AXI_NSV_M4
`endif 

`ifdef i_axi_AXI_LOG2_NSV_M4
  `define AXI_LOG2_NSV_M4 `i_axi_AXI_LOG2_NSV_M4
`endif 

`ifdef i_axi_AXI_NSV_M5
  `define AXI_NSV_M5 `i_axi_AXI_NSV_M5
`endif 

`ifdef i_axi_AXI_LOG2_NSV_M5
  `define AXI_LOG2_NSV_M5 `i_axi_AXI_LOG2_NSV_M5
`endif 

`ifdef i_axi_AXI_NSV_M6
  `define AXI_NSV_M6 `i_axi_AXI_NSV_M6
`endif 

`ifdef i_axi_AXI_LOG2_NSV_M6
  `define AXI_LOG2_NSV_M6 `i_axi_AXI_LOG2_NSV_M6
`endif 

`ifdef i_axi_AXI_NSV_M7
  `define AXI_NSV_M7 `i_axi_AXI_NSV_M7
`endif 

`ifdef i_axi_AXI_LOG2_NSV_M7
  `define AXI_LOG2_NSV_M7 `i_axi_AXI_LOG2_NSV_M7
`endif 

`ifdef i_axi_AXI_NSV_M8
  `define AXI_NSV_M8 `i_axi_AXI_NSV_M8
`endif 

`ifdef i_axi_AXI_LOG2_NSV_M8
  `define AXI_LOG2_NSV_M8 `i_axi_AXI_LOG2_NSV_M8
`endif 

`ifdef i_axi_AXI_NSV_M9
  `define AXI_NSV_M9 `i_axi_AXI_NSV_M9
`endif 

`ifdef i_axi_AXI_LOG2_NSV_M9
  `define AXI_LOG2_NSV_M9 `i_axi_AXI_LOG2_NSV_M9
`endif 

`ifdef i_axi_AXI_NSV_M10
  `define AXI_NSV_M10 `i_axi_AXI_NSV_M10
`endif 

`ifdef i_axi_AXI_LOG2_NSV_M10
  `define AXI_LOG2_NSV_M10 `i_axi_AXI_LOG2_NSV_M10
`endif 

`ifdef i_axi_AXI_NSV_M11
  `define AXI_NSV_M11 `i_axi_AXI_NSV_M11
`endif 

`ifdef i_axi_AXI_LOG2_NSV_M11
  `define AXI_LOG2_NSV_M11 `i_axi_AXI_LOG2_NSV_M11
`endif 

`ifdef i_axi_AXI_NSV_M12
  `define AXI_NSV_M12 `i_axi_AXI_NSV_M12
`endif 

`ifdef i_axi_AXI_LOG2_NSV_M12
  `define AXI_LOG2_NSV_M12 `i_axi_AXI_LOG2_NSV_M12
`endif 

`ifdef i_axi_AXI_NSV_M13
  `define AXI_NSV_M13 `i_axi_AXI_NSV_M13
`endif 

`ifdef i_axi_AXI_LOG2_NSV_M13
  `define AXI_LOG2_NSV_M13 `i_axi_AXI_LOG2_NSV_M13
`endif 

`ifdef i_axi_AXI_NSV_M14
  `define AXI_NSV_M14 `i_axi_AXI_NSV_M14
`endif 

`ifdef i_axi_AXI_LOG2_NSV_M14
  `define AXI_LOG2_NSV_M14 `i_axi_AXI_LOG2_NSV_M14
`endif 

`ifdef i_axi_AXI_NSV_M15
  `define AXI_NSV_M15 `i_axi_AXI_NSV_M15
`endif 

`ifdef i_axi_AXI_LOG2_NSV_M15
  `define AXI_LOG2_NSV_M15 `i_axi_AXI_LOG2_NSV_M15
`endif 

`ifdef i_axi_AXI_NSV_M16
  `define AXI_NSV_M16 `i_axi_AXI_NSV_M16
`endif 

`ifdef i_axi_AXI_LOG2_NSV_M16
  `define AXI_LOG2_NSV_M16 `i_axi_AXI_LOG2_NSV_M16
`endif 

`ifdef i_axi_AXI_NNMV_S1
  `define AXI_NNMV_S1 `i_axi_AXI_NNMV_S1
`endif 

`ifdef i_axi_AXI_BNMV_S1
  `define AXI_BNMV_S1 `i_axi_AXI_BNMV_S1
`endif 

`ifdef i_axi_AXI_NNMV_S2
  `define AXI_NNMV_S2 `i_axi_AXI_NNMV_S2
`endif 

`ifdef i_axi_AXI_BNMV_S2
  `define AXI_BNMV_S2 `i_axi_AXI_BNMV_S2
`endif 

`ifdef i_axi_AXI_NNMV_S3
  `define AXI_NNMV_S3 `i_axi_AXI_NNMV_S3
`endif 

`ifdef i_axi_AXI_BNMV_S3
  `define AXI_BNMV_S3 `i_axi_AXI_BNMV_S3
`endif 

`ifdef i_axi_AXI_NNMV_S4
  `define AXI_NNMV_S4 `i_axi_AXI_NNMV_S4
`endif 

`ifdef i_axi_AXI_BNMV_S4
  `define AXI_BNMV_S4 `i_axi_AXI_BNMV_S4
`endif 

`ifdef i_axi_AXI_NNMV_S5
  `define AXI_NNMV_S5 `i_axi_AXI_NNMV_S5
`endif 

`ifdef i_axi_AXI_BNMV_S5
  `define AXI_BNMV_S5 `i_axi_AXI_BNMV_S5
`endif 

`ifdef i_axi_AXI_NNMV_S6
  `define AXI_NNMV_S6 `i_axi_AXI_NNMV_S6
`endif 

`ifdef i_axi_AXI_BNMV_S6
  `define AXI_BNMV_S6 `i_axi_AXI_BNMV_S6
`endif 

`ifdef i_axi_AXI_NNMV_S7
  `define AXI_NNMV_S7 `i_axi_AXI_NNMV_S7
`endif 

`ifdef i_axi_AXI_BNMV_S7
  `define AXI_BNMV_S7 `i_axi_AXI_BNMV_S7
`endif 

`ifdef i_axi_AXI_NNMV_S8
  `define AXI_NNMV_S8 `i_axi_AXI_NNMV_S8
`endif 

`ifdef i_axi_AXI_BNMV_S8
  `define AXI_BNMV_S8 `i_axi_AXI_BNMV_S8
`endif 

`ifdef i_axi_AXI_NNMV_S9
  `define AXI_NNMV_S9 `i_axi_AXI_NNMV_S9
`endif 

`ifdef i_axi_AXI_BNMV_S9
  `define AXI_BNMV_S9 `i_axi_AXI_BNMV_S9
`endif 

`ifdef i_axi_AXI_NNMV_S10
  `define AXI_NNMV_S10 `i_axi_AXI_NNMV_S10
`endif 

`ifdef i_axi_AXI_BNMV_S10
  `define AXI_BNMV_S10 `i_axi_AXI_BNMV_S10
`endif 

`ifdef i_axi_AXI_NNMV_S11
  `define AXI_NNMV_S11 `i_axi_AXI_NNMV_S11
`endif 

`ifdef i_axi_AXI_BNMV_S11
  `define AXI_BNMV_S11 `i_axi_AXI_BNMV_S11
`endif 

`ifdef i_axi_AXI_NNMV_S12
  `define AXI_NNMV_S12 `i_axi_AXI_NNMV_S12
`endif 

`ifdef i_axi_AXI_BNMV_S12
  `define AXI_BNMV_S12 `i_axi_AXI_BNMV_S12
`endif 

`ifdef i_axi_AXI_NNMV_S13
  `define AXI_NNMV_S13 `i_axi_AXI_NNMV_S13
`endif 

`ifdef i_axi_AXI_BNMV_S13
  `define AXI_BNMV_S13 `i_axi_AXI_BNMV_S13
`endif 

`ifdef i_axi_AXI_NNMV_S14
  `define AXI_NNMV_S14 `i_axi_AXI_NNMV_S14
`endif 

`ifdef i_axi_AXI_BNMV_S14
  `define AXI_BNMV_S14 `i_axi_AXI_BNMV_S14
`endif 

`ifdef i_axi_AXI_NNMV_S15
  `define AXI_NNMV_S15 `i_axi_AXI_NNMV_S15
`endif 

`ifdef i_axi_AXI_BNMV_S15
  `define AXI_BNMV_S15 `i_axi_AXI_BNMV_S15
`endif 

`ifdef i_axi_AXI_NNMV_S16
  `define AXI_NNMV_S16 `i_axi_AXI_NNMV_S16
`endif 

`ifdef i_axi_AXI_BNMV_S16
  `define AXI_BNMV_S16 `i_axi_AXI_BNMV_S16
`endif 

`ifdef i_axi_AXI_NSP1V_M1
  `define AXI_NSP1V_M1 `i_axi_AXI_NSP1V_M1
`endif 

`ifdef i_axi_AXI_LOG2_NSP1V_M1
  `define AXI_LOG2_NSP1V_M1 `i_axi_AXI_LOG2_NSP1V_M1
`endif 

`ifdef i_axi_AXI_LOG2_NSP2V_M1
  `define AXI_LOG2_NSP2V_M1 `i_axi_AXI_LOG2_NSP2V_M1
`endif 

`ifdef i_axi_AXI_NSP1V_M2
  `define AXI_NSP1V_M2 `i_axi_AXI_NSP1V_M2
`endif 

`ifdef i_axi_AXI_LOG2_NSP1V_M2
  `define AXI_LOG2_NSP1V_M2 `i_axi_AXI_LOG2_NSP1V_M2
`endif 

`ifdef i_axi_AXI_LOG2_NSP2V_M2
  `define AXI_LOG2_NSP2V_M2 `i_axi_AXI_LOG2_NSP2V_M2
`endif 

`ifdef i_axi_AXI_NSP1V_M3
  `define AXI_NSP1V_M3 `i_axi_AXI_NSP1V_M3
`endif 

`ifdef i_axi_AXI_LOG2_NSP1V_M3
  `define AXI_LOG2_NSP1V_M3 `i_axi_AXI_LOG2_NSP1V_M3
`endif 

`ifdef i_axi_AXI_LOG2_NSP2V_M3
  `define AXI_LOG2_NSP2V_M3 `i_axi_AXI_LOG2_NSP2V_M3
`endif 

`ifdef i_axi_AXI_NSP1V_M4
  `define AXI_NSP1V_M4 `i_axi_AXI_NSP1V_M4
`endif 

`ifdef i_axi_AXI_LOG2_NSP1V_M4
  `define AXI_LOG2_NSP1V_M4 `i_axi_AXI_LOG2_NSP1V_M4
`endif 

`ifdef i_axi_AXI_LOG2_NSP2V_M4
  `define AXI_LOG2_NSP2V_M4 `i_axi_AXI_LOG2_NSP2V_M4
`endif 

`ifdef i_axi_AXI_NSP1V_M5
  `define AXI_NSP1V_M5 `i_axi_AXI_NSP1V_M5
`endif 

`ifdef i_axi_AXI_LOG2_NSP1V_M5
  `define AXI_LOG2_NSP1V_M5 `i_axi_AXI_LOG2_NSP1V_M5
`endif 

`ifdef i_axi_AXI_LOG2_NSP2V_M5
  `define AXI_LOG2_NSP2V_M5 `i_axi_AXI_LOG2_NSP2V_M5
`endif 

`ifdef i_axi_AXI_NSP1V_M6
  `define AXI_NSP1V_M6 `i_axi_AXI_NSP1V_M6
`endif 

`ifdef i_axi_AXI_LOG2_NSP1V_M6
  `define AXI_LOG2_NSP1V_M6 `i_axi_AXI_LOG2_NSP1V_M6
`endif 

`ifdef i_axi_AXI_LOG2_NSP2V_M6
  `define AXI_LOG2_NSP2V_M6 `i_axi_AXI_LOG2_NSP2V_M6
`endif 

`ifdef i_axi_AXI_NSP1V_M7
  `define AXI_NSP1V_M7 `i_axi_AXI_NSP1V_M7
`endif 

`ifdef i_axi_AXI_LOG2_NSP1V_M7
  `define AXI_LOG2_NSP1V_M7 `i_axi_AXI_LOG2_NSP1V_M7
`endif 

`ifdef i_axi_AXI_LOG2_NSP2V_M7
  `define AXI_LOG2_NSP2V_M7 `i_axi_AXI_LOG2_NSP2V_M7
`endif 

`ifdef i_axi_AXI_NSP1V_M8
  `define AXI_NSP1V_M8 `i_axi_AXI_NSP1V_M8
`endif 

`ifdef i_axi_AXI_LOG2_NSP1V_M8
  `define AXI_LOG2_NSP1V_M8 `i_axi_AXI_LOG2_NSP1V_M8
`endif 

`ifdef i_axi_AXI_LOG2_NSP2V_M8
  `define AXI_LOG2_NSP2V_M8 `i_axi_AXI_LOG2_NSP2V_M8
`endif 

`ifdef i_axi_AXI_NSP1V_M9
  `define AXI_NSP1V_M9 `i_axi_AXI_NSP1V_M9
`endif 

`ifdef i_axi_AXI_LOG2_NSP1V_M9
  `define AXI_LOG2_NSP1V_M9 `i_axi_AXI_LOG2_NSP1V_M9
`endif 

`ifdef i_axi_AXI_LOG2_NSP2V_M9
  `define AXI_LOG2_NSP2V_M9 `i_axi_AXI_LOG2_NSP2V_M9
`endif 

`ifdef i_axi_AXI_NSP1V_M10
  `define AXI_NSP1V_M10 `i_axi_AXI_NSP1V_M10
`endif 

`ifdef i_axi_AXI_LOG2_NSP1V_M10
  `define AXI_LOG2_NSP1V_M10 `i_axi_AXI_LOG2_NSP1V_M10
`endif 

`ifdef i_axi_AXI_LOG2_NSP2V_M10
  `define AXI_LOG2_NSP2V_M10 `i_axi_AXI_LOG2_NSP2V_M10
`endif 

`ifdef i_axi_AXI_NSP1V_M11
  `define AXI_NSP1V_M11 `i_axi_AXI_NSP1V_M11
`endif 

`ifdef i_axi_AXI_LOG2_NSP1V_M11
  `define AXI_LOG2_NSP1V_M11 `i_axi_AXI_LOG2_NSP1V_M11
`endif 

`ifdef i_axi_AXI_LOG2_NSP2V_M11
  `define AXI_LOG2_NSP2V_M11 `i_axi_AXI_LOG2_NSP2V_M11
`endif 

`ifdef i_axi_AXI_NSP1V_M12
  `define AXI_NSP1V_M12 `i_axi_AXI_NSP1V_M12
`endif 

`ifdef i_axi_AXI_LOG2_NSP1V_M12
  `define AXI_LOG2_NSP1V_M12 `i_axi_AXI_LOG2_NSP1V_M12
`endif 

`ifdef i_axi_AXI_LOG2_NSP2V_M12
  `define AXI_LOG2_NSP2V_M12 `i_axi_AXI_LOG2_NSP2V_M12
`endif 

`ifdef i_axi_AXI_NSP1V_M13
  `define AXI_NSP1V_M13 `i_axi_AXI_NSP1V_M13
`endif 

`ifdef i_axi_AXI_LOG2_NSP1V_M13
  `define AXI_LOG2_NSP1V_M13 `i_axi_AXI_LOG2_NSP1V_M13
`endif 

`ifdef i_axi_AXI_LOG2_NSP2V_M13
  `define AXI_LOG2_NSP2V_M13 `i_axi_AXI_LOG2_NSP2V_M13
`endif 

`ifdef i_axi_AXI_NSP1V_M14
  `define AXI_NSP1V_M14 `i_axi_AXI_NSP1V_M14
`endif 

`ifdef i_axi_AXI_LOG2_NSP1V_M14
  `define AXI_LOG2_NSP1V_M14 `i_axi_AXI_LOG2_NSP1V_M14
`endif 

`ifdef i_axi_AXI_LOG2_NSP2V_M14
  `define AXI_LOG2_NSP2V_M14 `i_axi_AXI_LOG2_NSP2V_M14
`endif 

`ifdef i_axi_AXI_NSP1V_M15
  `define AXI_NSP1V_M15 `i_axi_AXI_NSP1V_M15
`endif 

`ifdef i_axi_AXI_LOG2_NSP1V_M15
  `define AXI_LOG2_NSP1V_M15 `i_axi_AXI_LOG2_NSP1V_M15
`endif 

`ifdef i_axi_AXI_LOG2_NSP2V_M15
  `define AXI_LOG2_NSP2V_M15 `i_axi_AXI_LOG2_NSP2V_M15
`endif 

`ifdef i_axi_AXI_NSP1V_M16
  `define AXI_NSP1V_M16 `i_axi_AXI_NSP1V_M16
`endif 

`ifdef i_axi_AXI_LOG2_NSP1V_M16
  `define AXI_LOG2_NSP1V_M16 `i_axi_AXI_LOG2_NSP1V_M16
`endif 

`ifdef i_axi_AXI_LOG2_NSP2V_M16
  `define AXI_LOG2_NSP2V_M16 `i_axi_AXI_LOG2_NSP2V_M16
`endif 

`ifdef i_axi_AXI_ALL_AR_LAYER_SHARED
  `define AXI_ALL_AR_LAYER_SHARED `i_axi_AXI_ALL_AR_LAYER_SHARED
`endif 

`ifdef i_axi_AXI_AR_LAYER_S0_M1
  `define AXI_AR_LAYER_S0_M1 `i_axi_AXI_AR_LAYER_S0_M1
`endif 

`ifdef i_axi_AXI_AR_LAYER_S0_M2
  `define AXI_AR_LAYER_S0_M2 `i_axi_AXI_AR_LAYER_S0_M2
`endif 

`ifdef i_axi_AXI_AR_LAYER_S0_M3
  `define AXI_AR_LAYER_S0_M3 `i_axi_AXI_AR_LAYER_S0_M3
`endif 

`ifdef i_axi_AXI_AR_LAYER_S0_M4
  `define AXI_AR_LAYER_S0_M4 `i_axi_AXI_AR_LAYER_S0_M4
`endif 

`ifdef i_axi_AXI_AR_LAYER_S0_M5
  `define AXI_AR_LAYER_S0_M5 `i_axi_AXI_AR_LAYER_S0_M5
`endif 

`ifdef i_axi_AXI_AR_LAYER_S0_M6
  `define AXI_AR_LAYER_S0_M6 `i_axi_AXI_AR_LAYER_S0_M6
`endif 

`ifdef i_axi_AXI_AR_LAYER_S0_M7
  `define AXI_AR_LAYER_S0_M7 `i_axi_AXI_AR_LAYER_S0_M7
`endif 

`ifdef i_axi_AXI_AR_LAYER_S0_M8
  `define AXI_AR_LAYER_S0_M8 `i_axi_AXI_AR_LAYER_S0_M8
`endif 

`ifdef i_axi_AXI_AR_LAYER_S0_M9
  `define AXI_AR_LAYER_S0_M9 `i_axi_AXI_AR_LAYER_S0_M9
`endif 

`ifdef i_axi_AXI_AR_LAYER_S0_M10
  `define AXI_AR_LAYER_S0_M10 `i_axi_AXI_AR_LAYER_S0_M10
`endif 

`ifdef i_axi_AXI_AR_LAYER_S0_M11
  `define AXI_AR_LAYER_S0_M11 `i_axi_AXI_AR_LAYER_S0_M11
`endif 

`ifdef i_axi_AXI_AR_LAYER_S0_M12
  `define AXI_AR_LAYER_S0_M12 `i_axi_AXI_AR_LAYER_S0_M12
`endif 

`ifdef i_axi_AXI_AR_LAYER_S0_M13
  `define AXI_AR_LAYER_S0_M13 `i_axi_AXI_AR_LAYER_S0_M13
`endif 

`ifdef i_axi_AXI_AR_LAYER_S0_M14
  `define AXI_AR_LAYER_S0_M14 `i_axi_AXI_AR_LAYER_S0_M14
`endif 

`ifdef i_axi_AXI_AR_LAYER_S0_M15
  `define AXI_AR_LAYER_S0_M15 `i_axi_AXI_AR_LAYER_S0_M15
`endif 

`ifdef i_axi_AXI_AR_LAYER_S0_M16
  `define AXI_AR_LAYER_S0_M16 `i_axi_AXI_AR_LAYER_S0_M16
`endif 

`ifdef i_axi_AXI_ALL_AW_LAYER_SHARED
  `define AXI_ALL_AW_LAYER_SHARED `i_axi_AXI_ALL_AW_LAYER_SHARED
`endif 

`ifdef i_axi_AXI_AW_LAYER_S0_M1
  `define AXI_AW_LAYER_S0_M1 `i_axi_AXI_AW_LAYER_S0_M1
`endif 

`ifdef i_axi_AXI_AW_LAYER_S0_M2
  `define AXI_AW_LAYER_S0_M2 `i_axi_AXI_AW_LAYER_S0_M2
`endif 

`ifdef i_axi_AXI_AW_LAYER_S0_M3
  `define AXI_AW_LAYER_S0_M3 `i_axi_AXI_AW_LAYER_S0_M3
`endif 

`ifdef i_axi_AXI_AW_LAYER_S0_M4
  `define AXI_AW_LAYER_S0_M4 `i_axi_AXI_AW_LAYER_S0_M4
`endif 

`ifdef i_axi_AXI_AW_LAYER_S0_M5
  `define AXI_AW_LAYER_S0_M5 `i_axi_AXI_AW_LAYER_S0_M5
`endif 

`ifdef i_axi_AXI_AW_LAYER_S0_M6
  `define AXI_AW_LAYER_S0_M6 `i_axi_AXI_AW_LAYER_S0_M6
`endif 

`ifdef i_axi_AXI_AW_LAYER_S0_M7
  `define AXI_AW_LAYER_S0_M7 `i_axi_AXI_AW_LAYER_S0_M7
`endif 

`ifdef i_axi_AXI_AW_LAYER_S0_M8
  `define AXI_AW_LAYER_S0_M8 `i_axi_AXI_AW_LAYER_S0_M8
`endif 

`ifdef i_axi_AXI_AW_LAYER_S0_M9
  `define AXI_AW_LAYER_S0_M9 `i_axi_AXI_AW_LAYER_S0_M9
`endif 

`ifdef i_axi_AXI_AW_LAYER_S0_M10
  `define AXI_AW_LAYER_S0_M10 `i_axi_AXI_AW_LAYER_S0_M10
`endif 

`ifdef i_axi_AXI_AW_LAYER_S0_M11
  `define AXI_AW_LAYER_S0_M11 `i_axi_AXI_AW_LAYER_S0_M11
`endif 

`ifdef i_axi_AXI_AW_LAYER_S0_M12
  `define AXI_AW_LAYER_S0_M12 `i_axi_AXI_AW_LAYER_S0_M12
`endif 

`ifdef i_axi_AXI_AW_LAYER_S0_M13
  `define AXI_AW_LAYER_S0_M13 `i_axi_AXI_AW_LAYER_S0_M13
`endif 

`ifdef i_axi_AXI_AW_LAYER_S0_M14
  `define AXI_AW_LAYER_S0_M14 `i_axi_AXI_AW_LAYER_S0_M14
`endif 

`ifdef i_axi_AXI_AW_LAYER_S0_M15
  `define AXI_AW_LAYER_S0_M15 `i_axi_AXI_AW_LAYER_S0_M15
`endif 

`ifdef i_axi_AXI_AW_LAYER_S0_M16
  `define AXI_AW_LAYER_S0_M16 `i_axi_AXI_AW_LAYER_S0_M16
`endif 

`ifdef i_axi_AXI_ALL_W_LAYER_SHARED
  `define AXI_ALL_W_LAYER_SHARED `i_axi_AXI_ALL_W_LAYER_SHARED
`endif 

`ifdef i_axi_AXI_W_LAYER_S0_M1
  `define AXI_W_LAYER_S0_M1 `i_axi_AXI_W_LAYER_S0_M1
`endif 

`ifdef i_axi_AXI_W_LAYER_S0_M2
  `define AXI_W_LAYER_S0_M2 `i_axi_AXI_W_LAYER_S0_M2
`endif 

`ifdef i_axi_AXI_W_LAYER_S0_M3
  `define AXI_W_LAYER_S0_M3 `i_axi_AXI_W_LAYER_S0_M3
`endif 

`ifdef i_axi_AXI_W_LAYER_S0_M4
  `define AXI_W_LAYER_S0_M4 `i_axi_AXI_W_LAYER_S0_M4
`endif 

`ifdef i_axi_AXI_W_LAYER_S0_M5
  `define AXI_W_LAYER_S0_M5 `i_axi_AXI_W_LAYER_S0_M5
`endif 

`ifdef i_axi_AXI_W_LAYER_S0_M6
  `define AXI_W_LAYER_S0_M6 `i_axi_AXI_W_LAYER_S0_M6
`endif 

`ifdef i_axi_AXI_W_LAYER_S0_M7
  `define AXI_W_LAYER_S0_M7 `i_axi_AXI_W_LAYER_S0_M7
`endif 

`ifdef i_axi_AXI_W_LAYER_S0_M8
  `define AXI_W_LAYER_S0_M8 `i_axi_AXI_W_LAYER_S0_M8
`endif 

`ifdef i_axi_AXI_W_LAYER_S0_M9
  `define AXI_W_LAYER_S0_M9 `i_axi_AXI_W_LAYER_S0_M9
`endif 

`ifdef i_axi_AXI_W_LAYER_S0_M10
  `define AXI_W_LAYER_S0_M10 `i_axi_AXI_W_LAYER_S0_M10
`endif 

`ifdef i_axi_AXI_W_LAYER_S0_M11
  `define AXI_W_LAYER_S0_M11 `i_axi_AXI_W_LAYER_S0_M11
`endif 

`ifdef i_axi_AXI_W_LAYER_S0_M12
  `define AXI_W_LAYER_S0_M12 `i_axi_AXI_W_LAYER_S0_M12
`endif 

`ifdef i_axi_AXI_W_LAYER_S0_M13
  `define AXI_W_LAYER_S0_M13 `i_axi_AXI_W_LAYER_S0_M13
`endif 

`ifdef i_axi_AXI_W_LAYER_S0_M14
  `define AXI_W_LAYER_S0_M14 `i_axi_AXI_W_LAYER_S0_M14
`endif 

`ifdef i_axi_AXI_W_LAYER_S0_M15
  `define AXI_W_LAYER_S0_M15 `i_axi_AXI_W_LAYER_S0_M15
`endif 

`ifdef i_axi_AXI_W_LAYER_S0_M16
  `define AXI_W_LAYER_S0_M16 `i_axi_AXI_W_LAYER_S0_M16
`endif 

`ifdef i_axi_AXI_AR_LAYER_S1_M1
  `define AXI_AR_LAYER_S1_M1 `i_axi_AXI_AR_LAYER_S1_M1
`endif 

`ifdef i_axi_AXI_AR_LAYER_S1_M2
  `define AXI_AR_LAYER_S1_M2 `i_axi_AXI_AR_LAYER_S1_M2
`endif 

`ifdef i_axi_AXI_AR_LAYER_S1_M3
  `define AXI_AR_LAYER_S1_M3 `i_axi_AXI_AR_LAYER_S1_M3
`endif 

`ifdef i_axi_AXI_AR_LAYER_S1_M4
  `define AXI_AR_LAYER_S1_M4 `i_axi_AXI_AR_LAYER_S1_M4
`endif 

`ifdef i_axi_AXI_AR_LAYER_S1_M5
  `define AXI_AR_LAYER_S1_M5 `i_axi_AXI_AR_LAYER_S1_M5
`endif 

`ifdef i_axi_AXI_AR_LAYER_S1_M6
  `define AXI_AR_LAYER_S1_M6 `i_axi_AXI_AR_LAYER_S1_M6
`endif 

`ifdef i_axi_AXI_AR_LAYER_S1_M7
  `define AXI_AR_LAYER_S1_M7 `i_axi_AXI_AR_LAYER_S1_M7
`endif 

`ifdef i_axi_AXI_AR_LAYER_S1_M8
  `define AXI_AR_LAYER_S1_M8 `i_axi_AXI_AR_LAYER_S1_M8
`endif 

`ifdef i_axi_AXI_AR_LAYER_S1_M9
  `define AXI_AR_LAYER_S1_M9 `i_axi_AXI_AR_LAYER_S1_M9
`endif 

`ifdef i_axi_AXI_AR_LAYER_S1_M10
  `define AXI_AR_LAYER_S1_M10 `i_axi_AXI_AR_LAYER_S1_M10
`endif 

`ifdef i_axi_AXI_AR_LAYER_S1_M11
  `define AXI_AR_LAYER_S1_M11 `i_axi_AXI_AR_LAYER_S1_M11
`endif 

`ifdef i_axi_AXI_AR_LAYER_S1_M12
  `define AXI_AR_LAYER_S1_M12 `i_axi_AXI_AR_LAYER_S1_M12
`endif 

`ifdef i_axi_AXI_AR_LAYER_S1_M13
  `define AXI_AR_LAYER_S1_M13 `i_axi_AXI_AR_LAYER_S1_M13
`endif 

`ifdef i_axi_AXI_AR_LAYER_S1_M14
  `define AXI_AR_LAYER_S1_M14 `i_axi_AXI_AR_LAYER_S1_M14
`endif 

`ifdef i_axi_AXI_AR_LAYER_S1_M15
  `define AXI_AR_LAYER_S1_M15 `i_axi_AXI_AR_LAYER_S1_M15
`endif 

`ifdef i_axi_AXI_AR_LAYER_S1_M16
  `define AXI_AR_LAYER_S1_M16 `i_axi_AXI_AR_LAYER_S1_M16
`endif 

`ifdef i_axi_AXI_AW_LAYER_S1_M1
  `define AXI_AW_LAYER_S1_M1 `i_axi_AXI_AW_LAYER_S1_M1
`endif 

`ifdef i_axi_AXI_AW_LAYER_S1_M2
  `define AXI_AW_LAYER_S1_M2 `i_axi_AXI_AW_LAYER_S1_M2
`endif 

`ifdef i_axi_AXI_AW_LAYER_S1_M3
  `define AXI_AW_LAYER_S1_M3 `i_axi_AXI_AW_LAYER_S1_M3
`endif 

`ifdef i_axi_AXI_AW_LAYER_S1_M4
  `define AXI_AW_LAYER_S1_M4 `i_axi_AXI_AW_LAYER_S1_M4
`endif 

`ifdef i_axi_AXI_AW_LAYER_S1_M5
  `define AXI_AW_LAYER_S1_M5 `i_axi_AXI_AW_LAYER_S1_M5
`endif 

`ifdef i_axi_AXI_AW_LAYER_S1_M6
  `define AXI_AW_LAYER_S1_M6 `i_axi_AXI_AW_LAYER_S1_M6
`endif 

`ifdef i_axi_AXI_AW_LAYER_S1_M7
  `define AXI_AW_LAYER_S1_M7 `i_axi_AXI_AW_LAYER_S1_M7
`endif 

`ifdef i_axi_AXI_AW_LAYER_S1_M8
  `define AXI_AW_LAYER_S1_M8 `i_axi_AXI_AW_LAYER_S1_M8
`endif 

`ifdef i_axi_AXI_AW_LAYER_S1_M9
  `define AXI_AW_LAYER_S1_M9 `i_axi_AXI_AW_LAYER_S1_M9
`endif 

`ifdef i_axi_AXI_AW_LAYER_S1_M10
  `define AXI_AW_LAYER_S1_M10 `i_axi_AXI_AW_LAYER_S1_M10
`endif 

`ifdef i_axi_AXI_AW_LAYER_S1_M11
  `define AXI_AW_LAYER_S1_M11 `i_axi_AXI_AW_LAYER_S1_M11
`endif 

`ifdef i_axi_AXI_AW_LAYER_S1_M12
  `define AXI_AW_LAYER_S1_M12 `i_axi_AXI_AW_LAYER_S1_M12
`endif 

`ifdef i_axi_AXI_AW_LAYER_S1_M13
  `define AXI_AW_LAYER_S1_M13 `i_axi_AXI_AW_LAYER_S1_M13
`endif 

`ifdef i_axi_AXI_AW_LAYER_S1_M14
  `define AXI_AW_LAYER_S1_M14 `i_axi_AXI_AW_LAYER_S1_M14
`endif 

`ifdef i_axi_AXI_AW_LAYER_S1_M15
  `define AXI_AW_LAYER_S1_M15 `i_axi_AXI_AW_LAYER_S1_M15
`endif 

`ifdef i_axi_AXI_AW_LAYER_S1_M16
  `define AXI_AW_LAYER_S1_M16 `i_axi_AXI_AW_LAYER_S1_M16
`endif 

`ifdef i_axi_AXI_W_LAYER_S1_M1
  `define AXI_W_LAYER_S1_M1 `i_axi_AXI_W_LAYER_S1_M1
`endif 

`ifdef i_axi_AXI_W_LAYER_S1_M2
  `define AXI_W_LAYER_S1_M2 `i_axi_AXI_W_LAYER_S1_M2
`endif 

`ifdef i_axi_AXI_W_LAYER_S1_M3
  `define AXI_W_LAYER_S1_M3 `i_axi_AXI_W_LAYER_S1_M3
`endif 

`ifdef i_axi_AXI_W_LAYER_S1_M4
  `define AXI_W_LAYER_S1_M4 `i_axi_AXI_W_LAYER_S1_M4
`endif 

`ifdef i_axi_AXI_W_LAYER_S1_M5
  `define AXI_W_LAYER_S1_M5 `i_axi_AXI_W_LAYER_S1_M5
`endif 

`ifdef i_axi_AXI_W_LAYER_S1_M6
  `define AXI_W_LAYER_S1_M6 `i_axi_AXI_W_LAYER_S1_M6
`endif 

`ifdef i_axi_AXI_W_LAYER_S1_M7
  `define AXI_W_LAYER_S1_M7 `i_axi_AXI_W_LAYER_S1_M7
`endif 

`ifdef i_axi_AXI_W_LAYER_S1_M8
  `define AXI_W_LAYER_S1_M8 `i_axi_AXI_W_LAYER_S1_M8
`endif 

`ifdef i_axi_AXI_W_LAYER_S1_M9
  `define AXI_W_LAYER_S1_M9 `i_axi_AXI_W_LAYER_S1_M9
`endif 

`ifdef i_axi_AXI_W_LAYER_S1_M10
  `define AXI_W_LAYER_S1_M10 `i_axi_AXI_W_LAYER_S1_M10
`endif 

`ifdef i_axi_AXI_W_LAYER_S1_M11
  `define AXI_W_LAYER_S1_M11 `i_axi_AXI_W_LAYER_S1_M11
`endif 

`ifdef i_axi_AXI_W_LAYER_S1_M12
  `define AXI_W_LAYER_S1_M12 `i_axi_AXI_W_LAYER_S1_M12
`endif 

`ifdef i_axi_AXI_W_LAYER_S1_M13
  `define AXI_W_LAYER_S1_M13 `i_axi_AXI_W_LAYER_S1_M13
`endif 

`ifdef i_axi_AXI_W_LAYER_S1_M14
  `define AXI_W_LAYER_S1_M14 `i_axi_AXI_W_LAYER_S1_M14
`endif 

`ifdef i_axi_AXI_W_LAYER_S1_M15
  `define AXI_W_LAYER_S1_M15 `i_axi_AXI_W_LAYER_S1_M15
`endif 

`ifdef i_axi_AXI_W_LAYER_S1_M16
  `define AXI_W_LAYER_S1_M16 `i_axi_AXI_W_LAYER_S1_M16
`endif 

`ifdef i_axi_AXI_AR_LAYER_S2_M1
  `define AXI_AR_LAYER_S2_M1 `i_axi_AXI_AR_LAYER_S2_M1
`endif 

`ifdef i_axi_AXI_AR_LAYER_S2_M2
  `define AXI_AR_LAYER_S2_M2 `i_axi_AXI_AR_LAYER_S2_M2
`endif 

`ifdef i_axi_AXI_AR_LAYER_S2_M3
  `define AXI_AR_LAYER_S2_M3 `i_axi_AXI_AR_LAYER_S2_M3
`endif 

`ifdef i_axi_AXI_AR_LAYER_S2_M4
  `define AXI_AR_LAYER_S2_M4 `i_axi_AXI_AR_LAYER_S2_M4
`endif 

`ifdef i_axi_AXI_AR_LAYER_S2_M5
  `define AXI_AR_LAYER_S2_M5 `i_axi_AXI_AR_LAYER_S2_M5
`endif 

`ifdef i_axi_AXI_AR_LAYER_S2_M6
  `define AXI_AR_LAYER_S2_M6 `i_axi_AXI_AR_LAYER_S2_M6
`endif 

`ifdef i_axi_AXI_AR_LAYER_S2_M7
  `define AXI_AR_LAYER_S2_M7 `i_axi_AXI_AR_LAYER_S2_M7
`endif 

`ifdef i_axi_AXI_AR_LAYER_S2_M8
  `define AXI_AR_LAYER_S2_M8 `i_axi_AXI_AR_LAYER_S2_M8
`endif 

`ifdef i_axi_AXI_AR_LAYER_S2_M9
  `define AXI_AR_LAYER_S2_M9 `i_axi_AXI_AR_LAYER_S2_M9
`endif 

`ifdef i_axi_AXI_AR_LAYER_S2_M10
  `define AXI_AR_LAYER_S2_M10 `i_axi_AXI_AR_LAYER_S2_M10
`endif 

`ifdef i_axi_AXI_AR_LAYER_S2_M11
  `define AXI_AR_LAYER_S2_M11 `i_axi_AXI_AR_LAYER_S2_M11
`endif 

`ifdef i_axi_AXI_AR_LAYER_S2_M12
  `define AXI_AR_LAYER_S2_M12 `i_axi_AXI_AR_LAYER_S2_M12
`endif 

`ifdef i_axi_AXI_AR_LAYER_S2_M13
  `define AXI_AR_LAYER_S2_M13 `i_axi_AXI_AR_LAYER_S2_M13
`endif 

`ifdef i_axi_AXI_AR_LAYER_S2_M14
  `define AXI_AR_LAYER_S2_M14 `i_axi_AXI_AR_LAYER_S2_M14
`endif 

`ifdef i_axi_AXI_AR_LAYER_S2_M15
  `define AXI_AR_LAYER_S2_M15 `i_axi_AXI_AR_LAYER_S2_M15
`endif 

`ifdef i_axi_AXI_AR_LAYER_S2_M16
  `define AXI_AR_LAYER_S2_M16 `i_axi_AXI_AR_LAYER_S2_M16
`endif 

`ifdef i_axi_AXI_AW_LAYER_S2_M1
  `define AXI_AW_LAYER_S2_M1 `i_axi_AXI_AW_LAYER_S2_M1
`endif 

`ifdef i_axi_AXI_AW_LAYER_S2_M2
  `define AXI_AW_LAYER_S2_M2 `i_axi_AXI_AW_LAYER_S2_M2
`endif 

`ifdef i_axi_AXI_AW_LAYER_S2_M3
  `define AXI_AW_LAYER_S2_M3 `i_axi_AXI_AW_LAYER_S2_M3
`endif 

`ifdef i_axi_AXI_AW_LAYER_S2_M4
  `define AXI_AW_LAYER_S2_M4 `i_axi_AXI_AW_LAYER_S2_M4
`endif 

`ifdef i_axi_AXI_AW_LAYER_S2_M5
  `define AXI_AW_LAYER_S2_M5 `i_axi_AXI_AW_LAYER_S2_M5
`endif 

`ifdef i_axi_AXI_AW_LAYER_S2_M6
  `define AXI_AW_LAYER_S2_M6 `i_axi_AXI_AW_LAYER_S2_M6
`endif 

`ifdef i_axi_AXI_AW_LAYER_S2_M7
  `define AXI_AW_LAYER_S2_M7 `i_axi_AXI_AW_LAYER_S2_M7
`endif 

`ifdef i_axi_AXI_AW_LAYER_S2_M8
  `define AXI_AW_LAYER_S2_M8 `i_axi_AXI_AW_LAYER_S2_M8
`endif 

`ifdef i_axi_AXI_AW_LAYER_S2_M9
  `define AXI_AW_LAYER_S2_M9 `i_axi_AXI_AW_LAYER_S2_M9
`endif 

`ifdef i_axi_AXI_AW_LAYER_S2_M10
  `define AXI_AW_LAYER_S2_M10 `i_axi_AXI_AW_LAYER_S2_M10
`endif 

`ifdef i_axi_AXI_AW_LAYER_S2_M11
  `define AXI_AW_LAYER_S2_M11 `i_axi_AXI_AW_LAYER_S2_M11
`endif 

`ifdef i_axi_AXI_AW_LAYER_S2_M12
  `define AXI_AW_LAYER_S2_M12 `i_axi_AXI_AW_LAYER_S2_M12
`endif 

`ifdef i_axi_AXI_AW_LAYER_S2_M13
  `define AXI_AW_LAYER_S2_M13 `i_axi_AXI_AW_LAYER_S2_M13
`endif 

`ifdef i_axi_AXI_AW_LAYER_S2_M14
  `define AXI_AW_LAYER_S2_M14 `i_axi_AXI_AW_LAYER_S2_M14
`endif 

`ifdef i_axi_AXI_AW_LAYER_S2_M15
  `define AXI_AW_LAYER_S2_M15 `i_axi_AXI_AW_LAYER_S2_M15
`endif 

`ifdef i_axi_AXI_AW_LAYER_S2_M16
  `define AXI_AW_LAYER_S2_M16 `i_axi_AXI_AW_LAYER_S2_M16
`endif 

`ifdef i_axi_AXI_W_LAYER_S2_M1
  `define AXI_W_LAYER_S2_M1 `i_axi_AXI_W_LAYER_S2_M1
`endif 

`ifdef i_axi_AXI_W_LAYER_S2_M2
  `define AXI_W_LAYER_S2_M2 `i_axi_AXI_W_LAYER_S2_M2
`endif 

`ifdef i_axi_AXI_W_LAYER_S2_M3
  `define AXI_W_LAYER_S2_M3 `i_axi_AXI_W_LAYER_S2_M3
`endif 

`ifdef i_axi_AXI_W_LAYER_S2_M4
  `define AXI_W_LAYER_S2_M4 `i_axi_AXI_W_LAYER_S2_M4
`endif 

`ifdef i_axi_AXI_W_LAYER_S2_M5
  `define AXI_W_LAYER_S2_M5 `i_axi_AXI_W_LAYER_S2_M5
`endif 

`ifdef i_axi_AXI_W_LAYER_S2_M6
  `define AXI_W_LAYER_S2_M6 `i_axi_AXI_W_LAYER_S2_M6
`endif 

`ifdef i_axi_AXI_W_LAYER_S2_M7
  `define AXI_W_LAYER_S2_M7 `i_axi_AXI_W_LAYER_S2_M7
`endif 

`ifdef i_axi_AXI_W_LAYER_S2_M8
  `define AXI_W_LAYER_S2_M8 `i_axi_AXI_W_LAYER_S2_M8
`endif 

`ifdef i_axi_AXI_W_LAYER_S2_M9
  `define AXI_W_LAYER_S2_M9 `i_axi_AXI_W_LAYER_S2_M9
`endif 

`ifdef i_axi_AXI_W_LAYER_S2_M10
  `define AXI_W_LAYER_S2_M10 `i_axi_AXI_W_LAYER_S2_M10
`endif 

`ifdef i_axi_AXI_W_LAYER_S2_M11
  `define AXI_W_LAYER_S2_M11 `i_axi_AXI_W_LAYER_S2_M11
`endif 

`ifdef i_axi_AXI_W_LAYER_S2_M12
  `define AXI_W_LAYER_S2_M12 `i_axi_AXI_W_LAYER_S2_M12
`endif 

`ifdef i_axi_AXI_W_LAYER_S2_M13
  `define AXI_W_LAYER_S2_M13 `i_axi_AXI_W_LAYER_S2_M13
`endif 

`ifdef i_axi_AXI_W_LAYER_S2_M14
  `define AXI_W_LAYER_S2_M14 `i_axi_AXI_W_LAYER_S2_M14
`endif 

`ifdef i_axi_AXI_W_LAYER_S2_M15
  `define AXI_W_LAYER_S2_M15 `i_axi_AXI_W_LAYER_S2_M15
`endif 

`ifdef i_axi_AXI_W_LAYER_S2_M16
  `define AXI_W_LAYER_S2_M16 `i_axi_AXI_W_LAYER_S2_M16
`endif 

`ifdef i_axi_AXI_AR_LAYER_S3_M1
  `define AXI_AR_LAYER_S3_M1 `i_axi_AXI_AR_LAYER_S3_M1
`endif 

`ifdef i_axi_AXI_AR_LAYER_S3_M2
  `define AXI_AR_LAYER_S3_M2 `i_axi_AXI_AR_LAYER_S3_M2
`endif 

`ifdef i_axi_AXI_AR_LAYER_S3_M3
  `define AXI_AR_LAYER_S3_M3 `i_axi_AXI_AR_LAYER_S3_M3
`endif 

`ifdef i_axi_AXI_AR_LAYER_S3_M4
  `define AXI_AR_LAYER_S3_M4 `i_axi_AXI_AR_LAYER_S3_M4
`endif 

`ifdef i_axi_AXI_AR_LAYER_S3_M5
  `define AXI_AR_LAYER_S3_M5 `i_axi_AXI_AR_LAYER_S3_M5
`endif 

`ifdef i_axi_AXI_AR_LAYER_S3_M6
  `define AXI_AR_LAYER_S3_M6 `i_axi_AXI_AR_LAYER_S3_M6
`endif 

`ifdef i_axi_AXI_AR_LAYER_S3_M7
  `define AXI_AR_LAYER_S3_M7 `i_axi_AXI_AR_LAYER_S3_M7
`endif 

`ifdef i_axi_AXI_AR_LAYER_S3_M8
  `define AXI_AR_LAYER_S3_M8 `i_axi_AXI_AR_LAYER_S3_M8
`endif 

`ifdef i_axi_AXI_AR_LAYER_S3_M9
  `define AXI_AR_LAYER_S3_M9 `i_axi_AXI_AR_LAYER_S3_M9
`endif 

`ifdef i_axi_AXI_AR_LAYER_S3_M10
  `define AXI_AR_LAYER_S3_M10 `i_axi_AXI_AR_LAYER_S3_M10
`endif 

`ifdef i_axi_AXI_AR_LAYER_S3_M11
  `define AXI_AR_LAYER_S3_M11 `i_axi_AXI_AR_LAYER_S3_M11
`endif 

`ifdef i_axi_AXI_AR_LAYER_S3_M12
  `define AXI_AR_LAYER_S3_M12 `i_axi_AXI_AR_LAYER_S3_M12
`endif 

`ifdef i_axi_AXI_AR_LAYER_S3_M13
  `define AXI_AR_LAYER_S3_M13 `i_axi_AXI_AR_LAYER_S3_M13
`endif 

`ifdef i_axi_AXI_AR_LAYER_S3_M14
  `define AXI_AR_LAYER_S3_M14 `i_axi_AXI_AR_LAYER_S3_M14
`endif 

`ifdef i_axi_AXI_AR_LAYER_S3_M15
  `define AXI_AR_LAYER_S3_M15 `i_axi_AXI_AR_LAYER_S3_M15
`endif 

`ifdef i_axi_AXI_AR_LAYER_S3_M16
  `define AXI_AR_LAYER_S3_M16 `i_axi_AXI_AR_LAYER_S3_M16
`endif 

`ifdef i_axi_AXI_AW_LAYER_S3_M1
  `define AXI_AW_LAYER_S3_M1 `i_axi_AXI_AW_LAYER_S3_M1
`endif 

`ifdef i_axi_AXI_AW_LAYER_S3_M2
  `define AXI_AW_LAYER_S3_M2 `i_axi_AXI_AW_LAYER_S3_M2
`endif 

`ifdef i_axi_AXI_AW_LAYER_S3_M3
  `define AXI_AW_LAYER_S3_M3 `i_axi_AXI_AW_LAYER_S3_M3
`endif 

`ifdef i_axi_AXI_AW_LAYER_S3_M4
  `define AXI_AW_LAYER_S3_M4 `i_axi_AXI_AW_LAYER_S3_M4
`endif 

`ifdef i_axi_AXI_AW_LAYER_S3_M5
  `define AXI_AW_LAYER_S3_M5 `i_axi_AXI_AW_LAYER_S3_M5
`endif 

`ifdef i_axi_AXI_AW_LAYER_S3_M6
  `define AXI_AW_LAYER_S3_M6 `i_axi_AXI_AW_LAYER_S3_M6
`endif 

`ifdef i_axi_AXI_AW_LAYER_S3_M7
  `define AXI_AW_LAYER_S3_M7 `i_axi_AXI_AW_LAYER_S3_M7
`endif 

`ifdef i_axi_AXI_AW_LAYER_S3_M8
  `define AXI_AW_LAYER_S3_M8 `i_axi_AXI_AW_LAYER_S3_M8
`endif 

`ifdef i_axi_AXI_AW_LAYER_S3_M9
  `define AXI_AW_LAYER_S3_M9 `i_axi_AXI_AW_LAYER_S3_M9
`endif 

`ifdef i_axi_AXI_AW_LAYER_S3_M10
  `define AXI_AW_LAYER_S3_M10 `i_axi_AXI_AW_LAYER_S3_M10
`endif 

`ifdef i_axi_AXI_AW_LAYER_S3_M11
  `define AXI_AW_LAYER_S3_M11 `i_axi_AXI_AW_LAYER_S3_M11
`endif 

`ifdef i_axi_AXI_AW_LAYER_S3_M12
  `define AXI_AW_LAYER_S3_M12 `i_axi_AXI_AW_LAYER_S3_M12
`endif 

`ifdef i_axi_AXI_AW_LAYER_S3_M13
  `define AXI_AW_LAYER_S3_M13 `i_axi_AXI_AW_LAYER_S3_M13
`endif 

`ifdef i_axi_AXI_AW_LAYER_S3_M14
  `define AXI_AW_LAYER_S3_M14 `i_axi_AXI_AW_LAYER_S3_M14
`endif 

`ifdef i_axi_AXI_AW_LAYER_S3_M15
  `define AXI_AW_LAYER_S3_M15 `i_axi_AXI_AW_LAYER_S3_M15
`endif 

`ifdef i_axi_AXI_AW_LAYER_S3_M16
  `define AXI_AW_LAYER_S3_M16 `i_axi_AXI_AW_LAYER_S3_M16
`endif 

`ifdef i_axi_AXI_W_LAYER_S3_M1
  `define AXI_W_LAYER_S3_M1 `i_axi_AXI_W_LAYER_S3_M1
`endif 

`ifdef i_axi_AXI_W_LAYER_S3_M2
  `define AXI_W_LAYER_S3_M2 `i_axi_AXI_W_LAYER_S3_M2
`endif 

`ifdef i_axi_AXI_W_LAYER_S3_M3
  `define AXI_W_LAYER_S3_M3 `i_axi_AXI_W_LAYER_S3_M3
`endif 

`ifdef i_axi_AXI_W_LAYER_S3_M4
  `define AXI_W_LAYER_S3_M4 `i_axi_AXI_W_LAYER_S3_M4
`endif 

`ifdef i_axi_AXI_W_LAYER_S3_M5
  `define AXI_W_LAYER_S3_M5 `i_axi_AXI_W_LAYER_S3_M5
`endif 

`ifdef i_axi_AXI_W_LAYER_S3_M6
  `define AXI_W_LAYER_S3_M6 `i_axi_AXI_W_LAYER_S3_M6
`endif 

`ifdef i_axi_AXI_W_LAYER_S3_M7
  `define AXI_W_LAYER_S3_M7 `i_axi_AXI_W_LAYER_S3_M7
`endif 

`ifdef i_axi_AXI_W_LAYER_S3_M8
  `define AXI_W_LAYER_S3_M8 `i_axi_AXI_W_LAYER_S3_M8
`endif 

`ifdef i_axi_AXI_W_LAYER_S3_M9
  `define AXI_W_LAYER_S3_M9 `i_axi_AXI_W_LAYER_S3_M9
`endif 

`ifdef i_axi_AXI_W_LAYER_S3_M10
  `define AXI_W_LAYER_S3_M10 `i_axi_AXI_W_LAYER_S3_M10
`endif 

`ifdef i_axi_AXI_W_LAYER_S3_M11
  `define AXI_W_LAYER_S3_M11 `i_axi_AXI_W_LAYER_S3_M11
`endif 

`ifdef i_axi_AXI_W_LAYER_S3_M12
  `define AXI_W_LAYER_S3_M12 `i_axi_AXI_W_LAYER_S3_M12
`endif 

`ifdef i_axi_AXI_W_LAYER_S3_M13
  `define AXI_W_LAYER_S3_M13 `i_axi_AXI_W_LAYER_S3_M13
`endif 

`ifdef i_axi_AXI_W_LAYER_S3_M14
  `define AXI_W_LAYER_S3_M14 `i_axi_AXI_W_LAYER_S3_M14
`endif 

`ifdef i_axi_AXI_W_LAYER_S3_M15
  `define AXI_W_LAYER_S3_M15 `i_axi_AXI_W_LAYER_S3_M15
`endif 

`ifdef i_axi_AXI_W_LAYER_S3_M16
  `define AXI_W_LAYER_S3_M16 `i_axi_AXI_W_LAYER_S3_M16
`endif 

`ifdef i_axi_AXI_AR_LAYER_S4_M1
  `define AXI_AR_LAYER_S4_M1 `i_axi_AXI_AR_LAYER_S4_M1
`endif 

`ifdef i_axi_AXI_AR_LAYER_S4_M2
  `define AXI_AR_LAYER_S4_M2 `i_axi_AXI_AR_LAYER_S4_M2
`endif 

`ifdef i_axi_AXI_AR_LAYER_S4_M3
  `define AXI_AR_LAYER_S4_M3 `i_axi_AXI_AR_LAYER_S4_M3
`endif 

`ifdef i_axi_AXI_AR_LAYER_S4_M4
  `define AXI_AR_LAYER_S4_M4 `i_axi_AXI_AR_LAYER_S4_M4
`endif 

`ifdef i_axi_AXI_AR_LAYER_S4_M5
  `define AXI_AR_LAYER_S4_M5 `i_axi_AXI_AR_LAYER_S4_M5
`endif 

`ifdef i_axi_AXI_AR_LAYER_S4_M6
  `define AXI_AR_LAYER_S4_M6 `i_axi_AXI_AR_LAYER_S4_M6
`endif 

`ifdef i_axi_AXI_AR_LAYER_S4_M7
  `define AXI_AR_LAYER_S4_M7 `i_axi_AXI_AR_LAYER_S4_M7
`endif 

`ifdef i_axi_AXI_AR_LAYER_S4_M8
  `define AXI_AR_LAYER_S4_M8 `i_axi_AXI_AR_LAYER_S4_M8
`endif 

`ifdef i_axi_AXI_AR_LAYER_S4_M9
  `define AXI_AR_LAYER_S4_M9 `i_axi_AXI_AR_LAYER_S4_M9
`endif 

`ifdef i_axi_AXI_AR_LAYER_S4_M10
  `define AXI_AR_LAYER_S4_M10 `i_axi_AXI_AR_LAYER_S4_M10
`endif 

`ifdef i_axi_AXI_AR_LAYER_S4_M11
  `define AXI_AR_LAYER_S4_M11 `i_axi_AXI_AR_LAYER_S4_M11
`endif 

`ifdef i_axi_AXI_AR_LAYER_S4_M12
  `define AXI_AR_LAYER_S4_M12 `i_axi_AXI_AR_LAYER_S4_M12
`endif 

`ifdef i_axi_AXI_AR_LAYER_S4_M13
  `define AXI_AR_LAYER_S4_M13 `i_axi_AXI_AR_LAYER_S4_M13
`endif 

`ifdef i_axi_AXI_AR_LAYER_S4_M14
  `define AXI_AR_LAYER_S4_M14 `i_axi_AXI_AR_LAYER_S4_M14
`endif 

`ifdef i_axi_AXI_AR_LAYER_S4_M15
  `define AXI_AR_LAYER_S4_M15 `i_axi_AXI_AR_LAYER_S4_M15
`endif 

`ifdef i_axi_AXI_AR_LAYER_S4_M16
  `define AXI_AR_LAYER_S4_M16 `i_axi_AXI_AR_LAYER_S4_M16
`endif 

`ifdef i_axi_AXI_AW_LAYER_S4_M1
  `define AXI_AW_LAYER_S4_M1 `i_axi_AXI_AW_LAYER_S4_M1
`endif 

`ifdef i_axi_AXI_AW_LAYER_S4_M2
  `define AXI_AW_LAYER_S4_M2 `i_axi_AXI_AW_LAYER_S4_M2
`endif 

`ifdef i_axi_AXI_AW_LAYER_S4_M3
  `define AXI_AW_LAYER_S4_M3 `i_axi_AXI_AW_LAYER_S4_M3
`endif 

`ifdef i_axi_AXI_AW_LAYER_S4_M4
  `define AXI_AW_LAYER_S4_M4 `i_axi_AXI_AW_LAYER_S4_M4
`endif 

`ifdef i_axi_AXI_AW_LAYER_S4_M5
  `define AXI_AW_LAYER_S4_M5 `i_axi_AXI_AW_LAYER_S4_M5
`endif 

`ifdef i_axi_AXI_AW_LAYER_S4_M6
  `define AXI_AW_LAYER_S4_M6 `i_axi_AXI_AW_LAYER_S4_M6
`endif 

`ifdef i_axi_AXI_AW_LAYER_S4_M7
  `define AXI_AW_LAYER_S4_M7 `i_axi_AXI_AW_LAYER_S4_M7
`endif 

`ifdef i_axi_AXI_AW_LAYER_S4_M8
  `define AXI_AW_LAYER_S4_M8 `i_axi_AXI_AW_LAYER_S4_M8
`endif 

`ifdef i_axi_AXI_AW_LAYER_S4_M9
  `define AXI_AW_LAYER_S4_M9 `i_axi_AXI_AW_LAYER_S4_M9
`endif 

`ifdef i_axi_AXI_AW_LAYER_S4_M10
  `define AXI_AW_LAYER_S4_M10 `i_axi_AXI_AW_LAYER_S4_M10
`endif 

`ifdef i_axi_AXI_AW_LAYER_S4_M11
  `define AXI_AW_LAYER_S4_M11 `i_axi_AXI_AW_LAYER_S4_M11
`endif 

`ifdef i_axi_AXI_AW_LAYER_S4_M12
  `define AXI_AW_LAYER_S4_M12 `i_axi_AXI_AW_LAYER_S4_M12
`endif 

`ifdef i_axi_AXI_AW_LAYER_S4_M13
  `define AXI_AW_LAYER_S4_M13 `i_axi_AXI_AW_LAYER_S4_M13
`endif 

`ifdef i_axi_AXI_AW_LAYER_S4_M14
  `define AXI_AW_LAYER_S4_M14 `i_axi_AXI_AW_LAYER_S4_M14
`endif 

`ifdef i_axi_AXI_AW_LAYER_S4_M15
  `define AXI_AW_LAYER_S4_M15 `i_axi_AXI_AW_LAYER_S4_M15
`endif 

`ifdef i_axi_AXI_AW_LAYER_S4_M16
  `define AXI_AW_LAYER_S4_M16 `i_axi_AXI_AW_LAYER_S4_M16
`endif 

`ifdef i_axi_AXI_W_LAYER_S4_M1
  `define AXI_W_LAYER_S4_M1 `i_axi_AXI_W_LAYER_S4_M1
`endif 

`ifdef i_axi_AXI_W_LAYER_S4_M2
  `define AXI_W_LAYER_S4_M2 `i_axi_AXI_W_LAYER_S4_M2
`endif 

`ifdef i_axi_AXI_W_LAYER_S4_M3
  `define AXI_W_LAYER_S4_M3 `i_axi_AXI_W_LAYER_S4_M3
`endif 

`ifdef i_axi_AXI_W_LAYER_S4_M4
  `define AXI_W_LAYER_S4_M4 `i_axi_AXI_W_LAYER_S4_M4
`endif 

`ifdef i_axi_AXI_W_LAYER_S4_M5
  `define AXI_W_LAYER_S4_M5 `i_axi_AXI_W_LAYER_S4_M5
`endif 

`ifdef i_axi_AXI_W_LAYER_S4_M6
  `define AXI_W_LAYER_S4_M6 `i_axi_AXI_W_LAYER_S4_M6
`endif 

`ifdef i_axi_AXI_W_LAYER_S4_M7
  `define AXI_W_LAYER_S4_M7 `i_axi_AXI_W_LAYER_S4_M7
`endif 

`ifdef i_axi_AXI_W_LAYER_S4_M8
  `define AXI_W_LAYER_S4_M8 `i_axi_AXI_W_LAYER_S4_M8
`endif 

`ifdef i_axi_AXI_W_LAYER_S4_M9
  `define AXI_W_LAYER_S4_M9 `i_axi_AXI_W_LAYER_S4_M9
`endif 

`ifdef i_axi_AXI_W_LAYER_S4_M10
  `define AXI_W_LAYER_S4_M10 `i_axi_AXI_W_LAYER_S4_M10
`endif 

`ifdef i_axi_AXI_W_LAYER_S4_M11
  `define AXI_W_LAYER_S4_M11 `i_axi_AXI_W_LAYER_S4_M11
`endif 

`ifdef i_axi_AXI_W_LAYER_S4_M12
  `define AXI_W_LAYER_S4_M12 `i_axi_AXI_W_LAYER_S4_M12
`endif 

`ifdef i_axi_AXI_W_LAYER_S4_M13
  `define AXI_W_LAYER_S4_M13 `i_axi_AXI_W_LAYER_S4_M13
`endif 

`ifdef i_axi_AXI_W_LAYER_S4_M14
  `define AXI_W_LAYER_S4_M14 `i_axi_AXI_W_LAYER_S4_M14
`endif 

`ifdef i_axi_AXI_W_LAYER_S4_M15
  `define AXI_W_LAYER_S4_M15 `i_axi_AXI_W_LAYER_S4_M15
`endif 

`ifdef i_axi_AXI_W_LAYER_S4_M16
  `define AXI_W_LAYER_S4_M16 `i_axi_AXI_W_LAYER_S4_M16
`endif 

`ifdef i_axi_AXI_AR_LAYER_S5_M1
  `define AXI_AR_LAYER_S5_M1 `i_axi_AXI_AR_LAYER_S5_M1
`endif 

`ifdef i_axi_AXI_AR_LAYER_S5_M2
  `define AXI_AR_LAYER_S5_M2 `i_axi_AXI_AR_LAYER_S5_M2
`endif 

`ifdef i_axi_AXI_AR_LAYER_S5_M3
  `define AXI_AR_LAYER_S5_M3 `i_axi_AXI_AR_LAYER_S5_M3
`endif 

`ifdef i_axi_AXI_AR_LAYER_S5_M4
  `define AXI_AR_LAYER_S5_M4 `i_axi_AXI_AR_LAYER_S5_M4
`endif 

`ifdef i_axi_AXI_AR_LAYER_S5_M5
  `define AXI_AR_LAYER_S5_M5 `i_axi_AXI_AR_LAYER_S5_M5
`endif 

`ifdef i_axi_AXI_AR_LAYER_S5_M6
  `define AXI_AR_LAYER_S5_M6 `i_axi_AXI_AR_LAYER_S5_M6
`endif 

`ifdef i_axi_AXI_AR_LAYER_S5_M7
  `define AXI_AR_LAYER_S5_M7 `i_axi_AXI_AR_LAYER_S5_M7
`endif 

`ifdef i_axi_AXI_AR_LAYER_S5_M8
  `define AXI_AR_LAYER_S5_M8 `i_axi_AXI_AR_LAYER_S5_M8
`endif 

`ifdef i_axi_AXI_AR_LAYER_S5_M9
  `define AXI_AR_LAYER_S5_M9 `i_axi_AXI_AR_LAYER_S5_M9
`endif 

`ifdef i_axi_AXI_AR_LAYER_S5_M10
  `define AXI_AR_LAYER_S5_M10 `i_axi_AXI_AR_LAYER_S5_M10
`endif 

`ifdef i_axi_AXI_AR_LAYER_S5_M11
  `define AXI_AR_LAYER_S5_M11 `i_axi_AXI_AR_LAYER_S5_M11
`endif 

`ifdef i_axi_AXI_AR_LAYER_S5_M12
  `define AXI_AR_LAYER_S5_M12 `i_axi_AXI_AR_LAYER_S5_M12
`endif 

`ifdef i_axi_AXI_AR_LAYER_S5_M13
  `define AXI_AR_LAYER_S5_M13 `i_axi_AXI_AR_LAYER_S5_M13
`endif 

`ifdef i_axi_AXI_AR_LAYER_S5_M14
  `define AXI_AR_LAYER_S5_M14 `i_axi_AXI_AR_LAYER_S5_M14
`endif 

`ifdef i_axi_AXI_AR_LAYER_S5_M15
  `define AXI_AR_LAYER_S5_M15 `i_axi_AXI_AR_LAYER_S5_M15
`endif 

`ifdef i_axi_AXI_AR_LAYER_S5_M16
  `define AXI_AR_LAYER_S5_M16 `i_axi_AXI_AR_LAYER_S5_M16
`endif 

`ifdef i_axi_AXI_AW_LAYER_S5_M1
  `define AXI_AW_LAYER_S5_M1 `i_axi_AXI_AW_LAYER_S5_M1
`endif 

`ifdef i_axi_AXI_AW_LAYER_S5_M2
  `define AXI_AW_LAYER_S5_M2 `i_axi_AXI_AW_LAYER_S5_M2
`endif 

`ifdef i_axi_AXI_AW_LAYER_S5_M3
  `define AXI_AW_LAYER_S5_M3 `i_axi_AXI_AW_LAYER_S5_M3
`endif 

`ifdef i_axi_AXI_AW_LAYER_S5_M4
  `define AXI_AW_LAYER_S5_M4 `i_axi_AXI_AW_LAYER_S5_M4
`endif 

`ifdef i_axi_AXI_AW_LAYER_S5_M5
  `define AXI_AW_LAYER_S5_M5 `i_axi_AXI_AW_LAYER_S5_M5
`endif 

`ifdef i_axi_AXI_AW_LAYER_S5_M6
  `define AXI_AW_LAYER_S5_M6 `i_axi_AXI_AW_LAYER_S5_M6
`endif 

`ifdef i_axi_AXI_AW_LAYER_S5_M7
  `define AXI_AW_LAYER_S5_M7 `i_axi_AXI_AW_LAYER_S5_M7
`endif 

`ifdef i_axi_AXI_AW_LAYER_S5_M8
  `define AXI_AW_LAYER_S5_M8 `i_axi_AXI_AW_LAYER_S5_M8
`endif 

`ifdef i_axi_AXI_AW_LAYER_S5_M9
  `define AXI_AW_LAYER_S5_M9 `i_axi_AXI_AW_LAYER_S5_M9
`endif 

`ifdef i_axi_AXI_AW_LAYER_S5_M10
  `define AXI_AW_LAYER_S5_M10 `i_axi_AXI_AW_LAYER_S5_M10
`endif 

`ifdef i_axi_AXI_AW_LAYER_S5_M11
  `define AXI_AW_LAYER_S5_M11 `i_axi_AXI_AW_LAYER_S5_M11
`endif 

`ifdef i_axi_AXI_AW_LAYER_S5_M12
  `define AXI_AW_LAYER_S5_M12 `i_axi_AXI_AW_LAYER_S5_M12
`endif 

`ifdef i_axi_AXI_AW_LAYER_S5_M13
  `define AXI_AW_LAYER_S5_M13 `i_axi_AXI_AW_LAYER_S5_M13
`endif 

`ifdef i_axi_AXI_AW_LAYER_S5_M14
  `define AXI_AW_LAYER_S5_M14 `i_axi_AXI_AW_LAYER_S5_M14
`endif 

`ifdef i_axi_AXI_AW_LAYER_S5_M15
  `define AXI_AW_LAYER_S5_M15 `i_axi_AXI_AW_LAYER_S5_M15
`endif 

`ifdef i_axi_AXI_AW_LAYER_S5_M16
  `define AXI_AW_LAYER_S5_M16 `i_axi_AXI_AW_LAYER_S5_M16
`endif 

`ifdef i_axi_AXI_W_LAYER_S5_M1
  `define AXI_W_LAYER_S5_M1 `i_axi_AXI_W_LAYER_S5_M1
`endif 

`ifdef i_axi_AXI_W_LAYER_S5_M2
  `define AXI_W_LAYER_S5_M2 `i_axi_AXI_W_LAYER_S5_M2
`endif 

`ifdef i_axi_AXI_W_LAYER_S5_M3
  `define AXI_W_LAYER_S5_M3 `i_axi_AXI_W_LAYER_S5_M3
`endif 

`ifdef i_axi_AXI_W_LAYER_S5_M4
  `define AXI_W_LAYER_S5_M4 `i_axi_AXI_W_LAYER_S5_M4
`endif 

`ifdef i_axi_AXI_W_LAYER_S5_M5
  `define AXI_W_LAYER_S5_M5 `i_axi_AXI_W_LAYER_S5_M5
`endif 

`ifdef i_axi_AXI_W_LAYER_S5_M6
  `define AXI_W_LAYER_S5_M6 `i_axi_AXI_W_LAYER_S5_M6
`endif 

`ifdef i_axi_AXI_W_LAYER_S5_M7
  `define AXI_W_LAYER_S5_M7 `i_axi_AXI_W_LAYER_S5_M7
`endif 

`ifdef i_axi_AXI_W_LAYER_S5_M8
  `define AXI_W_LAYER_S5_M8 `i_axi_AXI_W_LAYER_S5_M8
`endif 

`ifdef i_axi_AXI_W_LAYER_S5_M9
  `define AXI_W_LAYER_S5_M9 `i_axi_AXI_W_LAYER_S5_M9
`endif 

`ifdef i_axi_AXI_W_LAYER_S5_M10
  `define AXI_W_LAYER_S5_M10 `i_axi_AXI_W_LAYER_S5_M10
`endif 

`ifdef i_axi_AXI_W_LAYER_S5_M11
  `define AXI_W_LAYER_S5_M11 `i_axi_AXI_W_LAYER_S5_M11
`endif 

`ifdef i_axi_AXI_W_LAYER_S5_M12
  `define AXI_W_LAYER_S5_M12 `i_axi_AXI_W_LAYER_S5_M12
`endif 

`ifdef i_axi_AXI_W_LAYER_S5_M13
  `define AXI_W_LAYER_S5_M13 `i_axi_AXI_W_LAYER_S5_M13
`endif 

`ifdef i_axi_AXI_W_LAYER_S5_M14
  `define AXI_W_LAYER_S5_M14 `i_axi_AXI_W_LAYER_S5_M14
`endif 

`ifdef i_axi_AXI_W_LAYER_S5_M15
  `define AXI_W_LAYER_S5_M15 `i_axi_AXI_W_LAYER_S5_M15
`endif 

`ifdef i_axi_AXI_W_LAYER_S5_M16
  `define AXI_W_LAYER_S5_M16 `i_axi_AXI_W_LAYER_S5_M16
`endif 

`ifdef i_axi_AXI_AR_LAYER_S6_M1
  `define AXI_AR_LAYER_S6_M1 `i_axi_AXI_AR_LAYER_S6_M1
`endif 

`ifdef i_axi_AXI_AR_LAYER_S6_M2
  `define AXI_AR_LAYER_S6_M2 `i_axi_AXI_AR_LAYER_S6_M2
`endif 

`ifdef i_axi_AXI_AR_LAYER_S6_M3
  `define AXI_AR_LAYER_S6_M3 `i_axi_AXI_AR_LAYER_S6_M3
`endif 

`ifdef i_axi_AXI_AR_LAYER_S6_M4
  `define AXI_AR_LAYER_S6_M4 `i_axi_AXI_AR_LAYER_S6_M4
`endif 

`ifdef i_axi_AXI_AR_LAYER_S6_M5
  `define AXI_AR_LAYER_S6_M5 `i_axi_AXI_AR_LAYER_S6_M5
`endif 

`ifdef i_axi_AXI_AR_LAYER_S6_M6
  `define AXI_AR_LAYER_S6_M6 `i_axi_AXI_AR_LAYER_S6_M6
`endif 

`ifdef i_axi_AXI_AR_LAYER_S6_M7
  `define AXI_AR_LAYER_S6_M7 `i_axi_AXI_AR_LAYER_S6_M7
`endif 

`ifdef i_axi_AXI_AR_LAYER_S6_M8
  `define AXI_AR_LAYER_S6_M8 `i_axi_AXI_AR_LAYER_S6_M8
`endif 

`ifdef i_axi_AXI_AR_LAYER_S6_M9
  `define AXI_AR_LAYER_S6_M9 `i_axi_AXI_AR_LAYER_S6_M9
`endif 

`ifdef i_axi_AXI_AR_LAYER_S6_M10
  `define AXI_AR_LAYER_S6_M10 `i_axi_AXI_AR_LAYER_S6_M10
`endif 

`ifdef i_axi_AXI_AR_LAYER_S6_M11
  `define AXI_AR_LAYER_S6_M11 `i_axi_AXI_AR_LAYER_S6_M11
`endif 

`ifdef i_axi_AXI_AR_LAYER_S6_M12
  `define AXI_AR_LAYER_S6_M12 `i_axi_AXI_AR_LAYER_S6_M12
`endif 

`ifdef i_axi_AXI_AR_LAYER_S6_M13
  `define AXI_AR_LAYER_S6_M13 `i_axi_AXI_AR_LAYER_S6_M13
`endif 

`ifdef i_axi_AXI_AR_LAYER_S6_M14
  `define AXI_AR_LAYER_S6_M14 `i_axi_AXI_AR_LAYER_S6_M14
`endif 

`ifdef i_axi_AXI_AR_LAYER_S6_M15
  `define AXI_AR_LAYER_S6_M15 `i_axi_AXI_AR_LAYER_S6_M15
`endif 

`ifdef i_axi_AXI_AR_LAYER_S6_M16
  `define AXI_AR_LAYER_S6_M16 `i_axi_AXI_AR_LAYER_S6_M16
`endif 

`ifdef i_axi_AXI_AW_LAYER_S6_M1
  `define AXI_AW_LAYER_S6_M1 `i_axi_AXI_AW_LAYER_S6_M1
`endif 

`ifdef i_axi_AXI_AW_LAYER_S6_M2
  `define AXI_AW_LAYER_S6_M2 `i_axi_AXI_AW_LAYER_S6_M2
`endif 

`ifdef i_axi_AXI_AW_LAYER_S6_M3
  `define AXI_AW_LAYER_S6_M3 `i_axi_AXI_AW_LAYER_S6_M3
`endif 

`ifdef i_axi_AXI_AW_LAYER_S6_M4
  `define AXI_AW_LAYER_S6_M4 `i_axi_AXI_AW_LAYER_S6_M4
`endif 

`ifdef i_axi_AXI_AW_LAYER_S6_M5
  `define AXI_AW_LAYER_S6_M5 `i_axi_AXI_AW_LAYER_S6_M5
`endif 

`ifdef i_axi_AXI_AW_LAYER_S6_M6
  `define AXI_AW_LAYER_S6_M6 `i_axi_AXI_AW_LAYER_S6_M6
`endif 

`ifdef i_axi_AXI_AW_LAYER_S6_M7
  `define AXI_AW_LAYER_S6_M7 `i_axi_AXI_AW_LAYER_S6_M7
`endif 

`ifdef i_axi_AXI_AW_LAYER_S6_M8
  `define AXI_AW_LAYER_S6_M8 `i_axi_AXI_AW_LAYER_S6_M8
`endif 

`ifdef i_axi_AXI_AW_LAYER_S6_M9
  `define AXI_AW_LAYER_S6_M9 `i_axi_AXI_AW_LAYER_S6_M9
`endif 

`ifdef i_axi_AXI_AW_LAYER_S6_M10
  `define AXI_AW_LAYER_S6_M10 `i_axi_AXI_AW_LAYER_S6_M10
`endif 

`ifdef i_axi_AXI_AW_LAYER_S6_M11
  `define AXI_AW_LAYER_S6_M11 `i_axi_AXI_AW_LAYER_S6_M11
`endif 

`ifdef i_axi_AXI_AW_LAYER_S6_M12
  `define AXI_AW_LAYER_S6_M12 `i_axi_AXI_AW_LAYER_S6_M12
`endif 

`ifdef i_axi_AXI_AW_LAYER_S6_M13
  `define AXI_AW_LAYER_S6_M13 `i_axi_AXI_AW_LAYER_S6_M13
`endif 

`ifdef i_axi_AXI_AW_LAYER_S6_M14
  `define AXI_AW_LAYER_S6_M14 `i_axi_AXI_AW_LAYER_S6_M14
`endif 

`ifdef i_axi_AXI_AW_LAYER_S6_M15
  `define AXI_AW_LAYER_S6_M15 `i_axi_AXI_AW_LAYER_S6_M15
`endif 

`ifdef i_axi_AXI_AW_LAYER_S6_M16
  `define AXI_AW_LAYER_S6_M16 `i_axi_AXI_AW_LAYER_S6_M16
`endif 

`ifdef i_axi_AXI_W_LAYER_S6_M1
  `define AXI_W_LAYER_S6_M1 `i_axi_AXI_W_LAYER_S6_M1
`endif 

`ifdef i_axi_AXI_W_LAYER_S6_M2
  `define AXI_W_LAYER_S6_M2 `i_axi_AXI_W_LAYER_S6_M2
`endif 

`ifdef i_axi_AXI_W_LAYER_S6_M3
  `define AXI_W_LAYER_S6_M3 `i_axi_AXI_W_LAYER_S6_M3
`endif 

`ifdef i_axi_AXI_W_LAYER_S6_M4
  `define AXI_W_LAYER_S6_M4 `i_axi_AXI_W_LAYER_S6_M4
`endif 

`ifdef i_axi_AXI_W_LAYER_S6_M5
  `define AXI_W_LAYER_S6_M5 `i_axi_AXI_W_LAYER_S6_M5
`endif 

`ifdef i_axi_AXI_W_LAYER_S6_M6
  `define AXI_W_LAYER_S6_M6 `i_axi_AXI_W_LAYER_S6_M6
`endif 

`ifdef i_axi_AXI_W_LAYER_S6_M7
  `define AXI_W_LAYER_S6_M7 `i_axi_AXI_W_LAYER_S6_M7
`endif 

`ifdef i_axi_AXI_W_LAYER_S6_M8
  `define AXI_W_LAYER_S6_M8 `i_axi_AXI_W_LAYER_S6_M8
`endif 

`ifdef i_axi_AXI_W_LAYER_S6_M9
  `define AXI_W_LAYER_S6_M9 `i_axi_AXI_W_LAYER_S6_M9
`endif 

`ifdef i_axi_AXI_W_LAYER_S6_M10
  `define AXI_W_LAYER_S6_M10 `i_axi_AXI_W_LAYER_S6_M10
`endif 

`ifdef i_axi_AXI_W_LAYER_S6_M11
  `define AXI_W_LAYER_S6_M11 `i_axi_AXI_W_LAYER_S6_M11
`endif 

`ifdef i_axi_AXI_W_LAYER_S6_M12
  `define AXI_W_LAYER_S6_M12 `i_axi_AXI_W_LAYER_S6_M12
`endif 

`ifdef i_axi_AXI_W_LAYER_S6_M13
  `define AXI_W_LAYER_S6_M13 `i_axi_AXI_W_LAYER_S6_M13
`endif 

`ifdef i_axi_AXI_W_LAYER_S6_M14
  `define AXI_W_LAYER_S6_M14 `i_axi_AXI_W_LAYER_S6_M14
`endif 

`ifdef i_axi_AXI_W_LAYER_S6_M15
  `define AXI_W_LAYER_S6_M15 `i_axi_AXI_W_LAYER_S6_M15
`endif 

`ifdef i_axi_AXI_W_LAYER_S6_M16
  `define AXI_W_LAYER_S6_M16 `i_axi_AXI_W_LAYER_S6_M16
`endif 

`ifdef i_axi_AXI_AR_LAYER_S7_M1
  `define AXI_AR_LAYER_S7_M1 `i_axi_AXI_AR_LAYER_S7_M1
`endif 

`ifdef i_axi_AXI_AR_LAYER_S7_M2
  `define AXI_AR_LAYER_S7_M2 `i_axi_AXI_AR_LAYER_S7_M2
`endif 

`ifdef i_axi_AXI_AR_LAYER_S7_M3
  `define AXI_AR_LAYER_S7_M3 `i_axi_AXI_AR_LAYER_S7_M3
`endif 

`ifdef i_axi_AXI_AR_LAYER_S7_M4
  `define AXI_AR_LAYER_S7_M4 `i_axi_AXI_AR_LAYER_S7_M4
`endif 

`ifdef i_axi_AXI_AR_LAYER_S7_M5
  `define AXI_AR_LAYER_S7_M5 `i_axi_AXI_AR_LAYER_S7_M5
`endif 

`ifdef i_axi_AXI_AR_LAYER_S7_M6
  `define AXI_AR_LAYER_S7_M6 `i_axi_AXI_AR_LAYER_S7_M6
`endif 

`ifdef i_axi_AXI_AR_LAYER_S7_M7
  `define AXI_AR_LAYER_S7_M7 `i_axi_AXI_AR_LAYER_S7_M7
`endif 

`ifdef i_axi_AXI_AR_LAYER_S7_M8
  `define AXI_AR_LAYER_S7_M8 `i_axi_AXI_AR_LAYER_S7_M8
`endif 

`ifdef i_axi_AXI_AR_LAYER_S7_M9
  `define AXI_AR_LAYER_S7_M9 `i_axi_AXI_AR_LAYER_S7_M9
`endif 

`ifdef i_axi_AXI_AR_LAYER_S7_M10
  `define AXI_AR_LAYER_S7_M10 `i_axi_AXI_AR_LAYER_S7_M10
`endif 

`ifdef i_axi_AXI_AR_LAYER_S7_M11
  `define AXI_AR_LAYER_S7_M11 `i_axi_AXI_AR_LAYER_S7_M11
`endif 

`ifdef i_axi_AXI_AR_LAYER_S7_M12
  `define AXI_AR_LAYER_S7_M12 `i_axi_AXI_AR_LAYER_S7_M12
`endif 

`ifdef i_axi_AXI_AR_LAYER_S7_M13
  `define AXI_AR_LAYER_S7_M13 `i_axi_AXI_AR_LAYER_S7_M13
`endif 

`ifdef i_axi_AXI_AR_LAYER_S7_M14
  `define AXI_AR_LAYER_S7_M14 `i_axi_AXI_AR_LAYER_S7_M14
`endif 

`ifdef i_axi_AXI_AR_LAYER_S7_M15
  `define AXI_AR_LAYER_S7_M15 `i_axi_AXI_AR_LAYER_S7_M15
`endif 

`ifdef i_axi_AXI_AR_LAYER_S7_M16
  `define AXI_AR_LAYER_S7_M16 `i_axi_AXI_AR_LAYER_S7_M16
`endif 

`ifdef i_axi_AXI_AW_LAYER_S7_M1
  `define AXI_AW_LAYER_S7_M1 `i_axi_AXI_AW_LAYER_S7_M1
`endif 

`ifdef i_axi_AXI_AW_LAYER_S7_M2
  `define AXI_AW_LAYER_S7_M2 `i_axi_AXI_AW_LAYER_S7_M2
`endif 

`ifdef i_axi_AXI_AW_LAYER_S7_M3
  `define AXI_AW_LAYER_S7_M3 `i_axi_AXI_AW_LAYER_S7_M3
`endif 

`ifdef i_axi_AXI_AW_LAYER_S7_M4
  `define AXI_AW_LAYER_S7_M4 `i_axi_AXI_AW_LAYER_S7_M4
`endif 

`ifdef i_axi_AXI_AW_LAYER_S7_M5
  `define AXI_AW_LAYER_S7_M5 `i_axi_AXI_AW_LAYER_S7_M5
`endif 

`ifdef i_axi_AXI_AW_LAYER_S7_M6
  `define AXI_AW_LAYER_S7_M6 `i_axi_AXI_AW_LAYER_S7_M6
`endif 

`ifdef i_axi_AXI_AW_LAYER_S7_M7
  `define AXI_AW_LAYER_S7_M7 `i_axi_AXI_AW_LAYER_S7_M7
`endif 

`ifdef i_axi_AXI_AW_LAYER_S7_M8
  `define AXI_AW_LAYER_S7_M8 `i_axi_AXI_AW_LAYER_S7_M8
`endif 

`ifdef i_axi_AXI_AW_LAYER_S7_M9
  `define AXI_AW_LAYER_S7_M9 `i_axi_AXI_AW_LAYER_S7_M9
`endif 

`ifdef i_axi_AXI_AW_LAYER_S7_M10
  `define AXI_AW_LAYER_S7_M10 `i_axi_AXI_AW_LAYER_S7_M10
`endif 

`ifdef i_axi_AXI_AW_LAYER_S7_M11
  `define AXI_AW_LAYER_S7_M11 `i_axi_AXI_AW_LAYER_S7_M11
`endif 

`ifdef i_axi_AXI_AW_LAYER_S7_M12
  `define AXI_AW_LAYER_S7_M12 `i_axi_AXI_AW_LAYER_S7_M12
`endif 

`ifdef i_axi_AXI_AW_LAYER_S7_M13
  `define AXI_AW_LAYER_S7_M13 `i_axi_AXI_AW_LAYER_S7_M13
`endif 

`ifdef i_axi_AXI_AW_LAYER_S7_M14
  `define AXI_AW_LAYER_S7_M14 `i_axi_AXI_AW_LAYER_S7_M14
`endif 

`ifdef i_axi_AXI_AW_LAYER_S7_M15
  `define AXI_AW_LAYER_S7_M15 `i_axi_AXI_AW_LAYER_S7_M15
`endif 

`ifdef i_axi_AXI_AW_LAYER_S7_M16
  `define AXI_AW_LAYER_S7_M16 `i_axi_AXI_AW_LAYER_S7_M16
`endif 

`ifdef i_axi_AXI_W_LAYER_S7_M1
  `define AXI_W_LAYER_S7_M1 `i_axi_AXI_W_LAYER_S7_M1
`endif 

`ifdef i_axi_AXI_W_LAYER_S7_M2
  `define AXI_W_LAYER_S7_M2 `i_axi_AXI_W_LAYER_S7_M2
`endif 

`ifdef i_axi_AXI_W_LAYER_S7_M3
  `define AXI_W_LAYER_S7_M3 `i_axi_AXI_W_LAYER_S7_M3
`endif 

`ifdef i_axi_AXI_W_LAYER_S7_M4
  `define AXI_W_LAYER_S7_M4 `i_axi_AXI_W_LAYER_S7_M4
`endif 

`ifdef i_axi_AXI_W_LAYER_S7_M5
  `define AXI_W_LAYER_S7_M5 `i_axi_AXI_W_LAYER_S7_M5
`endif 

`ifdef i_axi_AXI_W_LAYER_S7_M6
  `define AXI_W_LAYER_S7_M6 `i_axi_AXI_W_LAYER_S7_M6
`endif 

`ifdef i_axi_AXI_W_LAYER_S7_M7
  `define AXI_W_LAYER_S7_M7 `i_axi_AXI_W_LAYER_S7_M7
`endif 

`ifdef i_axi_AXI_W_LAYER_S7_M8
  `define AXI_W_LAYER_S7_M8 `i_axi_AXI_W_LAYER_S7_M8
`endif 

`ifdef i_axi_AXI_W_LAYER_S7_M9
  `define AXI_W_LAYER_S7_M9 `i_axi_AXI_W_LAYER_S7_M9
`endif 

`ifdef i_axi_AXI_W_LAYER_S7_M10
  `define AXI_W_LAYER_S7_M10 `i_axi_AXI_W_LAYER_S7_M10
`endif 

`ifdef i_axi_AXI_W_LAYER_S7_M11
  `define AXI_W_LAYER_S7_M11 `i_axi_AXI_W_LAYER_S7_M11
`endif 

`ifdef i_axi_AXI_W_LAYER_S7_M12
  `define AXI_W_LAYER_S7_M12 `i_axi_AXI_W_LAYER_S7_M12
`endif 

`ifdef i_axi_AXI_W_LAYER_S7_M13
  `define AXI_W_LAYER_S7_M13 `i_axi_AXI_W_LAYER_S7_M13
`endif 

`ifdef i_axi_AXI_W_LAYER_S7_M14
  `define AXI_W_LAYER_S7_M14 `i_axi_AXI_W_LAYER_S7_M14
`endif 

`ifdef i_axi_AXI_W_LAYER_S7_M15
  `define AXI_W_LAYER_S7_M15 `i_axi_AXI_W_LAYER_S7_M15
`endif 

`ifdef i_axi_AXI_W_LAYER_S7_M16
  `define AXI_W_LAYER_S7_M16 `i_axi_AXI_W_LAYER_S7_M16
`endif 

`ifdef i_axi_AXI_AR_LAYER_S8_M1
  `define AXI_AR_LAYER_S8_M1 `i_axi_AXI_AR_LAYER_S8_M1
`endif 

`ifdef i_axi_AXI_AR_LAYER_S8_M2
  `define AXI_AR_LAYER_S8_M2 `i_axi_AXI_AR_LAYER_S8_M2
`endif 

`ifdef i_axi_AXI_AR_LAYER_S8_M3
  `define AXI_AR_LAYER_S8_M3 `i_axi_AXI_AR_LAYER_S8_M3
`endif 

`ifdef i_axi_AXI_AR_LAYER_S8_M4
  `define AXI_AR_LAYER_S8_M4 `i_axi_AXI_AR_LAYER_S8_M4
`endif 

`ifdef i_axi_AXI_AR_LAYER_S8_M5
  `define AXI_AR_LAYER_S8_M5 `i_axi_AXI_AR_LAYER_S8_M5
`endif 

`ifdef i_axi_AXI_AR_LAYER_S8_M6
  `define AXI_AR_LAYER_S8_M6 `i_axi_AXI_AR_LAYER_S8_M6
`endif 

`ifdef i_axi_AXI_AR_LAYER_S8_M7
  `define AXI_AR_LAYER_S8_M7 `i_axi_AXI_AR_LAYER_S8_M7
`endif 

`ifdef i_axi_AXI_AR_LAYER_S8_M8
  `define AXI_AR_LAYER_S8_M8 `i_axi_AXI_AR_LAYER_S8_M8
`endif 

`ifdef i_axi_AXI_AR_LAYER_S8_M9
  `define AXI_AR_LAYER_S8_M9 `i_axi_AXI_AR_LAYER_S8_M9
`endif 

`ifdef i_axi_AXI_AR_LAYER_S8_M10
  `define AXI_AR_LAYER_S8_M10 `i_axi_AXI_AR_LAYER_S8_M10
`endif 

`ifdef i_axi_AXI_AR_LAYER_S8_M11
  `define AXI_AR_LAYER_S8_M11 `i_axi_AXI_AR_LAYER_S8_M11
`endif 

`ifdef i_axi_AXI_AR_LAYER_S8_M12
  `define AXI_AR_LAYER_S8_M12 `i_axi_AXI_AR_LAYER_S8_M12
`endif 

`ifdef i_axi_AXI_AR_LAYER_S8_M13
  `define AXI_AR_LAYER_S8_M13 `i_axi_AXI_AR_LAYER_S8_M13
`endif 

`ifdef i_axi_AXI_AR_LAYER_S8_M14
  `define AXI_AR_LAYER_S8_M14 `i_axi_AXI_AR_LAYER_S8_M14
`endif 

`ifdef i_axi_AXI_AR_LAYER_S8_M15
  `define AXI_AR_LAYER_S8_M15 `i_axi_AXI_AR_LAYER_S8_M15
`endif 

`ifdef i_axi_AXI_AR_LAYER_S8_M16
  `define AXI_AR_LAYER_S8_M16 `i_axi_AXI_AR_LAYER_S8_M16
`endif 

`ifdef i_axi_AXI_AW_LAYER_S8_M1
  `define AXI_AW_LAYER_S8_M1 `i_axi_AXI_AW_LAYER_S8_M1
`endif 

`ifdef i_axi_AXI_AW_LAYER_S8_M2
  `define AXI_AW_LAYER_S8_M2 `i_axi_AXI_AW_LAYER_S8_M2
`endif 

`ifdef i_axi_AXI_AW_LAYER_S8_M3
  `define AXI_AW_LAYER_S8_M3 `i_axi_AXI_AW_LAYER_S8_M3
`endif 

`ifdef i_axi_AXI_AW_LAYER_S8_M4
  `define AXI_AW_LAYER_S8_M4 `i_axi_AXI_AW_LAYER_S8_M4
`endif 

`ifdef i_axi_AXI_AW_LAYER_S8_M5
  `define AXI_AW_LAYER_S8_M5 `i_axi_AXI_AW_LAYER_S8_M5
`endif 

`ifdef i_axi_AXI_AW_LAYER_S8_M6
  `define AXI_AW_LAYER_S8_M6 `i_axi_AXI_AW_LAYER_S8_M6
`endif 

`ifdef i_axi_AXI_AW_LAYER_S8_M7
  `define AXI_AW_LAYER_S8_M7 `i_axi_AXI_AW_LAYER_S8_M7
`endif 

`ifdef i_axi_AXI_AW_LAYER_S8_M8
  `define AXI_AW_LAYER_S8_M8 `i_axi_AXI_AW_LAYER_S8_M8
`endif 

`ifdef i_axi_AXI_AW_LAYER_S8_M9
  `define AXI_AW_LAYER_S8_M9 `i_axi_AXI_AW_LAYER_S8_M9
`endif 

`ifdef i_axi_AXI_AW_LAYER_S8_M10
  `define AXI_AW_LAYER_S8_M10 `i_axi_AXI_AW_LAYER_S8_M10
`endif 

`ifdef i_axi_AXI_AW_LAYER_S8_M11
  `define AXI_AW_LAYER_S8_M11 `i_axi_AXI_AW_LAYER_S8_M11
`endif 

`ifdef i_axi_AXI_AW_LAYER_S8_M12
  `define AXI_AW_LAYER_S8_M12 `i_axi_AXI_AW_LAYER_S8_M12
`endif 

`ifdef i_axi_AXI_AW_LAYER_S8_M13
  `define AXI_AW_LAYER_S8_M13 `i_axi_AXI_AW_LAYER_S8_M13
`endif 

`ifdef i_axi_AXI_AW_LAYER_S8_M14
  `define AXI_AW_LAYER_S8_M14 `i_axi_AXI_AW_LAYER_S8_M14
`endif 

`ifdef i_axi_AXI_AW_LAYER_S8_M15
  `define AXI_AW_LAYER_S8_M15 `i_axi_AXI_AW_LAYER_S8_M15
`endif 

`ifdef i_axi_AXI_AW_LAYER_S8_M16
  `define AXI_AW_LAYER_S8_M16 `i_axi_AXI_AW_LAYER_S8_M16
`endif 

`ifdef i_axi_AXI_W_LAYER_S8_M1
  `define AXI_W_LAYER_S8_M1 `i_axi_AXI_W_LAYER_S8_M1
`endif 

`ifdef i_axi_AXI_W_LAYER_S8_M2
  `define AXI_W_LAYER_S8_M2 `i_axi_AXI_W_LAYER_S8_M2
`endif 

`ifdef i_axi_AXI_W_LAYER_S8_M3
  `define AXI_W_LAYER_S8_M3 `i_axi_AXI_W_LAYER_S8_M3
`endif 

`ifdef i_axi_AXI_W_LAYER_S8_M4
  `define AXI_W_LAYER_S8_M4 `i_axi_AXI_W_LAYER_S8_M4
`endif 

`ifdef i_axi_AXI_W_LAYER_S8_M5
  `define AXI_W_LAYER_S8_M5 `i_axi_AXI_W_LAYER_S8_M5
`endif 

`ifdef i_axi_AXI_W_LAYER_S8_M6
  `define AXI_W_LAYER_S8_M6 `i_axi_AXI_W_LAYER_S8_M6
`endif 

`ifdef i_axi_AXI_W_LAYER_S8_M7
  `define AXI_W_LAYER_S8_M7 `i_axi_AXI_W_LAYER_S8_M7
`endif 

`ifdef i_axi_AXI_W_LAYER_S8_M8
  `define AXI_W_LAYER_S8_M8 `i_axi_AXI_W_LAYER_S8_M8
`endif 

`ifdef i_axi_AXI_W_LAYER_S8_M9
  `define AXI_W_LAYER_S8_M9 `i_axi_AXI_W_LAYER_S8_M9
`endif 

`ifdef i_axi_AXI_W_LAYER_S8_M10
  `define AXI_W_LAYER_S8_M10 `i_axi_AXI_W_LAYER_S8_M10
`endif 

`ifdef i_axi_AXI_W_LAYER_S8_M11
  `define AXI_W_LAYER_S8_M11 `i_axi_AXI_W_LAYER_S8_M11
`endif 

`ifdef i_axi_AXI_W_LAYER_S8_M12
  `define AXI_W_LAYER_S8_M12 `i_axi_AXI_W_LAYER_S8_M12
`endif 

`ifdef i_axi_AXI_W_LAYER_S8_M13
  `define AXI_W_LAYER_S8_M13 `i_axi_AXI_W_LAYER_S8_M13
`endif 

`ifdef i_axi_AXI_W_LAYER_S8_M14
  `define AXI_W_LAYER_S8_M14 `i_axi_AXI_W_LAYER_S8_M14
`endif 

`ifdef i_axi_AXI_W_LAYER_S8_M15
  `define AXI_W_LAYER_S8_M15 `i_axi_AXI_W_LAYER_S8_M15
`endif 

`ifdef i_axi_AXI_W_LAYER_S8_M16
  `define AXI_W_LAYER_S8_M16 `i_axi_AXI_W_LAYER_S8_M16
`endif 

`ifdef i_axi_AXI_AR_LAYER_S9_M1
  `define AXI_AR_LAYER_S9_M1 `i_axi_AXI_AR_LAYER_S9_M1
`endif 

`ifdef i_axi_AXI_AR_LAYER_S9_M2
  `define AXI_AR_LAYER_S9_M2 `i_axi_AXI_AR_LAYER_S9_M2
`endif 

`ifdef i_axi_AXI_AR_LAYER_S9_M3
  `define AXI_AR_LAYER_S9_M3 `i_axi_AXI_AR_LAYER_S9_M3
`endif 

`ifdef i_axi_AXI_AR_LAYER_S9_M4
  `define AXI_AR_LAYER_S9_M4 `i_axi_AXI_AR_LAYER_S9_M4
`endif 

`ifdef i_axi_AXI_AR_LAYER_S9_M5
  `define AXI_AR_LAYER_S9_M5 `i_axi_AXI_AR_LAYER_S9_M5
`endif 

`ifdef i_axi_AXI_AR_LAYER_S9_M6
  `define AXI_AR_LAYER_S9_M6 `i_axi_AXI_AR_LAYER_S9_M6
`endif 

`ifdef i_axi_AXI_AR_LAYER_S9_M7
  `define AXI_AR_LAYER_S9_M7 `i_axi_AXI_AR_LAYER_S9_M7
`endif 

`ifdef i_axi_AXI_AR_LAYER_S9_M8
  `define AXI_AR_LAYER_S9_M8 `i_axi_AXI_AR_LAYER_S9_M8
`endif 

`ifdef i_axi_AXI_AR_LAYER_S9_M9
  `define AXI_AR_LAYER_S9_M9 `i_axi_AXI_AR_LAYER_S9_M9
`endif 

`ifdef i_axi_AXI_AR_LAYER_S9_M10
  `define AXI_AR_LAYER_S9_M10 `i_axi_AXI_AR_LAYER_S9_M10
`endif 

`ifdef i_axi_AXI_AR_LAYER_S9_M11
  `define AXI_AR_LAYER_S9_M11 `i_axi_AXI_AR_LAYER_S9_M11
`endif 

`ifdef i_axi_AXI_AR_LAYER_S9_M12
  `define AXI_AR_LAYER_S9_M12 `i_axi_AXI_AR_LAYER_S9_M12
`endif 

`ifdef i_axi_AXI_AR_LAYER_S9_M13
  `define AXI_AR_LAYER_S9_M13 `i_axi_AXI_AR_LAYER_S9_M13
`endif 

`ifdef i_axi_AXI_AR_LAYER_S9_M14
  `define AXI_AR_LAYER_S9_M14 `i_axi_AXI_AR_LAYER_S9_M14
`endif 

`ifdef i_axi_AXI_AR_LAYER_S9_M15
  `define AXI_AR_LAYER_S9_M15 `i_axi_AXI_AR_LAYER_S9_M15
`endif 

`ifdef i_axi_AXI_AR_LAYER_S9_M16
  `define AXI_AR_LAYER_S9_M16 `i_axi_AXI_AR_LAYER_S9_M16
`endif 

`ifdef i_axi_AXI_AW_LAYER_S9_M1
  `define AXI_AW_LAYER_S9_M1 `i_axi_AXI_AW_LAYER_S9_M1
`endif 

`ifdef i_axi_AXI_AW_LAYER_S9_M2
  `define AXI_AW_LAYER_S9_M2 `i_axi_AXI_AW_LAYER_S9_M2
`endif 

`ifdef i_axi_AXI_AW_LAYER_S9_M3
  `define AXI_AW_LAYER_S9_M3 `i_axi_AXI_AW_LAYER_S9_M3
`endif 

`ifdef i_axi_AXI_AW_LAYER_S9_M4
  `define AXI_AW_LAYER_S9_M4 `i_axi_AXI_AW_LAYER_S9_M4
`endif 

`ifdef i_axi_AXI_AW_LAYER_S9_M5
  `define AXI_AW_LAYER_S9_M5 `i_axi_AXI_AW_LAYER_S9_M5
`endif 

`ifdef i_axi_AXI_AW_LAYER_S9_M6
  `define AXI_AW_LAYER_S9_M6 `i_axi_AXI_AW_LAYER_S9_M6
`endif 

`ifdef i_axi_AXI_AW_LAYER_S9_M7
  `define AXI_AW_LAYER_S9_M7 `i_axi_AXI_AW_LAYER_S9_M7
`endif 

`ifdef i_axi_AXI_AW_LAYER_S9_M8
  `define AXI_AW_LAYER_S9_M8 `i_axi_AXI_AW_LAYER_S9_M8
`endif 

`ifdef i_axi_AXI_AW_LAYER_S9_M9
  `define AXI_AW_LAYER_S9_M9 `i_axi_AXI_AW_LAYER_S9_M9
`endif 

`ifdef i_axi_AXI_AW_LAYER_S9_M10
  `define AXI_AW_LAYER_S9_M10 `i_axi_AXI_AW_LAYER_S9_M10
`endif 

`ifdef i_axi_AXI_AW_LAYER_S9_M11
  `define AXI_AW_LAYER_S9_M11 `i_axi_AXI_AW_LAYER_S9_M11
`endif 

`ifdef i_axi_AXI_AW_LAYER_S9_M12
  `define AXI_AW_LAYER_S9_M12 `i_axi_AXI_AW_LAYER_S9_M12
`endif 

`ifdef i_axi_AXI_AW_LAYER_S9_M13
  `define AXI_AW_LAYER_S9_M13 `i_axi_AXI_AW_LAYER_S9_M13
`endif 

`ifdef i_axi_AXI_AW_LAYER_S9_M14
  `define AXI_AW_LAYER_S9_M14 `i_axi_AXI_AW_LAYER_S9_M14
`endif 

`ifdef i_axi_AXI_AW_LAYER_S9_M15
  `define AXI_AW_LAYER_S9_M15 `i_axi_AXI_AW_LAYER_S9_M15
`endif 

`ifdef i_axi_AXI_AW_LAYER_S9_M16
  `define AXI_AW_LAYER_S9_M16 `i_axi_AXI_AW_LAYER_S9_M16
`endif 

`ifdef i_axi_AXI_W_LAYER_S9_M1
  `define AXI_W_LAYER_S9_M1 `i_axi_AXI_W_LAYER_S9_M1
`endif 

`ifdef i_axi_AXI_W_LAYER_S9_M2
  `define AXI_W_LAYER_S9_M2 `i_axi_AXI_W_LAYER_S9_M2
`endif 

`ifdef i_axi_AXI_W_LAYER_S9_M3
  `define AXI_W_LAYER_S9_M3 `i_axi_AXI_W_LAYER_S9_M3
`endif 

`ifdef i_axi_AXI_W_LAYER_S9_M4
  `define AXI_W_LAYER_S9_M4 `i_axi_AXI_W_LAYER_S9_M4
`endif 

`ifdef i_axi_AXI_W_LAYER_S9_M5
  `define AXI_W_LAYER_S9_M5 `i_axi_AXI_W_LAYER_S9_M5
`endif 

`ifdef i_axi_AXI_W_LAYER_S9_M6
  `define AXI_W_LAYER_S9_M6 `i_axi_AXI_W_LAYER_S9_M6
`endif 

`ifdef i_axi_AXI_W_LAYER_S9_M7
  `define AXI_W_LAYER_S9_M7 `i_axi_AXI_W_LAYER_S9_M7
`endif 

`ifdef i_axi_AXI_W_LAYER_S9_M8
  `define AXI_W_LAYER_S9_M8 `i_axi_AXI_W_LAYER_S9_M8
`endif 

`ifdef i_axi_AXI_W_LAYER_S9_M9
  `define AXI_W_LAYER_S9_M9 `i_axi_AXI_W_LAYER_S9_M9
`endif 

`ifdef i_axi_AXI_W_LAYER_S9_M10
  `define AXI_W_LAYER_S9_M10 `i_axi_AXI_W_LAYER_S9_M10
`endif 

`ifdef i_axi_AXI_W_LAYER_S9_M11
  `define AXI_W_LAYER_S9_M11 `i_axi_AXI_W_LAYER_S9_M11
`endif 

`ifdef i_axi_AXI_W_LAYER_S9_M12
  `define AXI_W_LAYER_S9_M12 `i_axi_AXI_W_LAYER_S9_M12
`endif 

`ifdef i_axi_AXI_W_LAYER_S9_M13
  `define AXI_W_LAYER_S9_M13 `i_axi_AXI_W_LAYER_S9_M13
`endif 

`ifdef i_axi_AXI_W_LAYER_S9_M14
  `define AXI_W_LAYER_S9_M14 `i_axi_AXI_W_LAYER_S9_M14
`endif 

`ifdef i_axi_AXI_W_LAYER_S9_M15
  `define AXI_W_LAYER_S9_M15 `i_axi_AXI_W_LAYER_S9_M15
`endif 

`ifdef i_axi_AXI_W_LAYER_S9_M16
  `define AXI_W_LAYER_S9_M16 `i_axi_AXI_W_LAYER_S9_M16
`endif 

`ifdef i_axi_AXI_AR_LAYER_S10_M1
  `define AXI_AR_LAYER_S10_M1 `i_axi_AXI_AR_LAYER_S10_M1
`endif 

`ifdef i_axi_AXI_AR_LAYER_S10_M2
  `define AXI_AR_LAYER_S10_M2 `i_axi_AXI_AR_LAYER_S10_M2
`endif 

`ifdef i_axi_AXI_AR_LAYER_S10_M3
  `define AXI_AR_LAYER_S10_M3 `i_axi_AXI_AR_LAYER_S10_M3
`endif 

`ifdef i_axi_AXI_AR_LAYER_S10_M4
  `define AXI_AR_LAYER_S10_M4 `i_axi_AXI_AR_LAYER_S10_M4
`endif 

`ifdef i_axi_AXI_AR_LAYER_S10_M5
  `define AXI_AR_LAYER_S10_M5 `i_axi_AXI_AR_LAYER_S10_M5
`endif 

`ifdef i_axi_AXI_AR_LAYER_S10_M6
  `define AXI_AR_LAYER_S10_M6 `i_axi_AXI_AR_LAYER_S10_M6
`endif 

`ifdef i_axi_AXI_AR_LAYER_S10_M7
  `define AXI_AR_LAYER_S10_M7 `i_axi_AXI_AR_LAYER_S10_M7
`endif 

`ifdef i_axi_AXI_AR_LAYER_S10_M8
  `define AXI_AR_LAYER_S10_M8 `i_axi_AXI_AR_LAYER_S10_M8
`endif 

`ifdef i_axi_AXI_AR_LAYER_S10_M9
  `define AXI_AR_LAYER_S10_M9 `i_axi_AXI_AR_LAYER_S10_M9
`endif 

`ifdef i_axi_AXI_AR_LAYER_S10_M10
  `define AXI_AR_LAYER_S10_M10 `i_axi_AXI_AR_LAYER_S10_M10
`endif 

`ifdef i_axi_AXI_AR_LAYER_S10_M11
  `define AXI_AR_LAYER_S10_M11 `i_axi_AXI_AR_LAYER_S10_M11
`endif 

`ifdef i_axi_AXI_AR_LAYER_S10_M12
  `define AXI_AR_LAYER_S10_M12 `i_axi_AXI_AR_LAYER_S10_M12
`endif 

`ifdef i_axi_AXI_AR_LAYER_S10_M13
  `define AXI_AR_LAYER_S10_M13 `i_axi_AXI_AR_LAYER_S10_M13
`endif 

`ifdef i_axi_AXI_AR_LAYER_S10_M14
  `define AXI_AR_LAYER_S10_M14 `i_axi_AXI_AR_LAYER_S10_M14
`endif 

`ifdef i_axi_AXI_AR_LAYER_S10_M15
  `define AXI_AR_LAYER_S10_M15 `i_axi_AXI_AR_LAYER_S10_M15
`endif 

`ifdef i_axi_AXI_AR_LAYER_S10_M16
  `define AXI_AR_LAYER_S10_M16 `i_axi_AXI_AR_LAYER_S10_M16
`endif 

`ifdef i_axi_AXI_AW_LAYER_S10_M1
  `define AXI_AW_LAYER_S10_M1 `i_axi_AXI_AW_LAYER_S10_M1
`endif 

`ifdef i_axi_AXI_AW_LAYER_S10_M2
  `define AXI_AW_LAYER_S10_M2 `i_axi_AXI_AW_LAYER_S10_M2
`endif 

`ifdef i_axi_AXI_AW_LAYER_S10_M3
  `define AXI_AW_LAYER_S10_M3 `i_axi_AXI_AW_LAYER_S10_M3
`endif 

`ifdef i_axi_AXI_AW_LAYER_S10_M4
  `define AXI_AW_LAYER_S10_M4 `i_axi_AXI_AW_LAYER_S10_M4
`endif 

`ifdef i_axi_AXI_AW_LAYER_S10_M5
  `define AXI_AW_LAYER_S10_M5 `i_axi_AXI_AW_LAYER_S10_M5
`endif 

`ifdef i_axi_AXI_AW_LAYER_S10_M6
  `define AXI_AW_LAYER_S10_M6 `i_axi_AXI_AW_LAYER_S10_M6
`endif 

`ifdef i_axi_AXI_AW_LAYER_S10_M7
  `define AXI_AW_LAYER_S10_M7 `i_axi_AXI_AW_LAYER_S10_M7
`endif 

`ifdef i_axi_AXI_AW_LAYER_S10_M8
  `define AXI_AW_LAYER_S10_M8 `i_axi_AXI_AW_LAYER_S10_M8
`endif 

`ifdef i_axi_AXI_AW_LAYER_S10_M9
  `define AXI_AW_LAYER_S10_M9 `i_axi_AXI_AW_LAYER_S10_M9
`endif 

`ifdef i_axi_AXI_AW_LAYER_S10_M10
  `define AXI_AW_LAYER_S10_M10 `i_axi_AXI_AW_LAYER_S10_M10
`endif 

`ifdef i_axi_AXI_AW_LAYER_S10_M11
  `define AXI_AW_LAYER_S10_M11 `i_axi_AXI_AW_LAYER_S10_M11
`endif 

`ifdef i_axi_AXI_AW_LAYER_S10_M12
  `define AXI_AW_LAYER_S10_M12 `i_axi_AXI_AW_LAYER_S10_M12
`endif 

`ifdef i_axi_AXI_AW_LAYER_S10_M13
  `define AXI_AW_LAYER_S10_M13 `i_axi_AXI_AW_LAYER_S10_M13
`endif 

`ifdef i_axi_AXI_AW_LAYER_S10_M14
  `define AXI_AW_LAYER_S10_M14 `i_axi_AXI_AW_LAYER_S10_M14
`endif 

`ifdef i_axi_AXI_AW_LAYER_S10_M15
  `define AXI_AW_LAYER_S10_M15 `i_axi_AXI_AW_LAYER_S10_M15
`endif 

`ifdef i_axi_AXI_AW_LAYER_S10_M16
  `define AXI_AW_LAYER_S10_M16 `i_axi_AXI_AW_LAYER_S10_M16
`endif 

`ifdef i_axi_AXI_W_LAYER_S10_M1
  `define AXI_W_LAYER_S10_M1 `i_axi_AXI_W_LAYER_S10_M1
`endif 

`ifdef i_axi_AXI_W_LAYER_S10_M2
  `define AXI_W_LAYER_S10_M2 `i_axi_AXI_W_LAYER_S10_M2
`endif 

`ifdef i_axi_AXI_W_LAYER_S10_M3
  `define AXI_W_LAYER_S10_M3 `i_axi_AXI_W_LAYER_S10_M3
`endif 

`ifdef i_axi_AXI_W_LAYER_S10_M4
  `define AXI_W_LAYER_S10_M4 `i_axi_AXI_W_LAYER_S10_M4
`endif 

`ifdef i_axi_AXI_W_LAYER_S10_M5
  `define AXI_W_LAYER_S10_M5 `i_axi_AXI_W_LAYER_S10_M5
`endif 

`ifdef i_axi_AXI_W_LAYER_S10_M6
  `define AXI_W_LAYER_S10_M6 `i_axi_AXI_W_LAYER_S10_M6
`endif 

`ifdef i_axi_AXI_W_LAYER_S10_M7
  `define AXI_W_LAYER_S10_M7 `i_axi_AXI_W_LAYER_S10_M7
`endif 

`ifdef i_axi_AXI_W_LAYER_S10_M8
  `define AXI_W_LAYER_S10_M8 `i_axi_AXI_W_LAYER_S10_M8
`endif 

`ifdef i_axi_AXI_W_LAYER_S10_M9
  `define AXI_W_LAYER_S10_M9 `i_axi_AXI_W_LAYER_S10_M9
`endif 

`ifdef i_axi_AXI_W_LAYER_S10_M10
  `define AXI_W_LAYER_S10_M10 `i_axi_AXI_W_LAYER_S10_M10
`endif 

`ifdef i_axi_AXI_W_LAYER_S10_M11
  `define AXI_W_LAYER_S10_M11 `i_axi_AXI_W_LAYER_S10_M11
`endif 

`ifdef i_axi_AXI_W_LAYER_S10_M12
  `define AXI_W_LAYER_S10_M12 `i_axi_AXI_W_LAYER_S10_M12
`endif 

`ifdef i_axi_AXI_W_LAYER_S10_M13
  `define AXI_W_LAYER_S10_M13 `i_axi_AXI_W_LAYER_S10_M13
`endif 

`ifdef i_axi_AXI_W_LAYER_S10_M14
  `define AXI_W_LAYER_S10_M14 `i_axi_AXI_W_LAYER_S10_M14
`endif 

`ifdef i_axi_AXI_W_LAYER_S10_M15
  `define AXI_W_LAYER_S10_M15 `i_axi_AXI_W_LAYER_S10_M15
`endif 

`ifdef i_axi_AXI_W_LAYER_S10_M16
  `define AXI_W_LAYER_S10_M16 `i_axi_AXI_W_LAYER_S10_M16
`endif 

`ifdef i_axi_AXI_AR_LAYER_S11_M1
  `define AXI_AR_LAYER_S11_M1 `i_axi_AXI_AR_LAYER_S11_M1
`endif 

`ifdef i_axi_AXI_AR_LAYER_S11_M2
  `define AXI_AR_LAYER_S11_M2 `i_axi_AXI_AR_LAYER_S11_M2
`endif 

`ifdef i_axi_AXI_AR_LAYER_S11_M3
  `define AXI_AR_LAYER_S11_M3 `i_axi_AXI_AR_LAYER_S11_M3
`endif 

`ifdef i_axi_AXI_AR_LAYER_S11_M4
  `define AXI_AR_LAYER_S11_M4 `i_axi_AXI_AR_LAYER_S11_M4
`endif 

`ifdef i_axi_AXI_AR_LAYER_S11_M5
  `define AXI_AR_LAYER_S11_M5 `i_axi_AXI_AR_LAYER_S11_M5
`endif 

`ifdef i_axi_AXI_AR_LAYER_S11_M6
  `define AXI_AR_LAYER_S11_M6 `i_axi_AXI_AR_LAYER_S11_M6
`endif 

`ifdef i_axi_AXI_AR_LAYER_S11_M7
  `define AXI_AR_LAYER_S11_M7 `i_axi_AXI_AR_LAYER_S11_M7
`endif 

`ifdef i_axi_AXI_AR_LAYER_S11_M8
  `define AXI_AR_LAYER_S11_M8 `i_axi_AXI_AR_LAYER_S11_M8
`endif 

`ifdef i_axi_AXI_AR_LAYER_S11_M9
  `define AXI_AR_LAYER_S11_M9 `i_axi_AXI_AR_LAYER_S11_M9
`endif 

`ifdef i_axi_AXI_AR_LAYER_S11_M10
  `define AXI_AR_LAYER_S11_M10 `i_axi_AXI_AR_LAYER_S11_M10
`endif 

`ifdef i_axi_AXI_AR_LAYER_S11_M11
  `define AXI_AR_LAYER_S11_M11 `i_axi_AXI_AR_LAYER_S11_M11
`endif 

`ifdef i_axi_AXI_AR_LAYER_S11_M12
  `define AXI_AR_LAYER_S11_M12 `i_axi_AXI_AR_LAYER_S11_M12
`endif 

`ifdef i_axi_AXI_AR_LAYER_S11_M13
  `define AXI_AR_LAYER_S11_M13 `i_axi_AXI_AR_LAYER_S11_M13
`endif 

`ifdef i_axi_AXI_AR_LAYER_S11_M14
  `define AXI_AR_LAYER_S11_M14 `i_axi_AXI_AR_LAYER_S11_M14
`endif 

`ifdef i_axi_AXI_AR_LAYER_S11_M15
  `define AXI_AR_LAYER_S11_M15 `i_axi_AXI_AR_LAYER_S11_M15
`endif 

`ifdef i_axi_AXI_AR_LAYER_S11_M16
  `define AXI_AR_LAYER_S11_M16 `i_axi_AXI_AR_LAYER_S11_M16
`endif 

`ifdef i_axi_AXI_AW_LAYER_S11_M1
  `define AXI_AW_LAYER_S11_M1 `i_axi_AXI_AW_LAYER_S11_M1
`endif 

`ifdef i_axi_AXI_AW_LAYER_S11_M2
  `define AXI_AW_LAYER_S11_M2 `i_axi_AXI_AW_LAYER_S11_M2
`endif 

`ifdef i_axi_AXI_AW_LAYER_S11_M3
  `define AXI_AW_LAYER_S11_M3 `i_axi_AXI_AW_LAYER_S11_M3
`endif 

`ifdef i_axi_AXI_AW_LAYER_S11_M4
  `define AXI_AW_LAYER_S11_M4 `i_axi_AXI_AW_LAYER_S11_M4
`endif 

`ifdef i_axi_AXI_AW_LAYER_S11_M5
  `define AXI_AW_LAYER_S11_M5 `i_axi_AXI_AW_LAYER_S11_M5
`endif 

`ifdef i_axi_AXI_AW_LAYER_S11_M6
  `define AXI_AW_LAYER_S11_M6 `i_axi_AXI_AW_LAYER_S11_M6
`endif 

`ifdef i_axi_AXI_AW_LAYER_S11_M7
  `define AXI_AW_LAYER_S11_M7 `i_axi_AXI_AW_LAYER_S11_M7
`endif 

`ifdef i_axi_AXI_AW_LAYER_S11_M8
  `define AXI_AW_LAYER_S11_M8 `i_axi_AXI_AW_LAYER_S11_M8
`endif 

`ifdef i_axi_AXI_AW_LAYER_S11_M9
  `define AXI_AW_LAYER_S11_M9 `i_axi_AXI_AW_LAYER_S11_M9
`endif 

`ifdef i_axi_AXI_AW_LAYER_S11_M10
  `define AXI_AW_LAYER_S11_M10 `i_axi_AXI_AW_LAYER_S11_M10
`endif 

`ifdef i_axi_AXI_AW_LAYER_S11_M11
  `define AXI_AW_LAYER_S11_M11 `i_axi_AXI_AW_LAYER_S11_M11
`endif 

`ifdef i_axi_AXI_AW_LAYER_S11_M12
  `define AXI_AW_LAYER_S11_M12 `i_axi_AXI_AW_LAYER_S11_M12
`endif 

`ifdef i_axi_AXI_AW_LAYER_S11_M13
  `define AXI_AW_LAYER_S11_M13 `i_axi_AXI_AW_LAYER_S11_M13
`endif 

`ifdef i_axi_AXI_AW_LAYER_S11_M14
  `define AXI_AW_LAYER_S11_M14 `i_axi_AXI_AW_LAYER_S11_M14
`endif 

`ifdef i_axi_AXI_AW_LAYER_S11_M15
  `define AXI_AW_LAYER_S11_M15 `i_axi_AXI_AW_LAYER_S11_M15
`endif 

`ifdef i_axi_AXI_AW_LAYER_S11_M16
  `define AXI_AW_LAYER_S11_M16 `i_axi_AXI_AW_LAYER_S11_M16
`endif 

`ifdef i_axi_AXI_W_LAYER_S11_M1
  `define AXI_W_LAYER_S11_M1 `i_axi_AXI_W_LAYER_S11_M1
`endif 

`ifdef i_axi_AXI_W_LAYER_S11_M2
  `define AXI_W_LAYER_S11_M2 `i_axi_AXI_W_LAYER_S11_M2
`endif 

`ifdef i_axi_AXI_W_LAYER_S11_M3
  `define AXI_W_LAYER_S11_M3 `i_axi_AXI_W_LAYER_S11_M3
`endif 

`ifdef i_axi_AXI_W_LAYER_S11_M4
  `define AXI_W_LAYER_S11_M4 `i_axi_AXI_W_LAYER_S11_M4
`endif 

`ifdef i_axi_AXI_W_LAYER_S11_M5
  `define AXI_W_LAYER_S11_M5 `i_axi_AXI_W_LAYER_S11_M5
`endif 

`ifdef i_axi_AXI_W_LAYER_S11_M6
  `define AXI_W_LAYER_S11_M6 `i_axi_AXI_W_LAYER_S11_M6
`endif 

`ifdef i_axi_AXI_W_LAYER_S11_M7
  `define AXI_W_LAYER_S11_M7 `i_axi_AXI_W_LAYER_S11_M7
`endif 

`ifdef i_axi_AXI_W_LAYER_S11_M8
  `define AXI_W_LAYER_S11_M8 `i_axi_AXI_W_LAYER_S11_M8
`endif 

`ifdef i_axi_AXI_W_LAYER_S11_M9
  `define AXI_W_LAYER_S11_M9 `i_axi_AXI_W_LAYER_S11_M9
`endif 

`ifdef i_axi_AXI_W_LAYER_S11_M10
  `define AXI_W_LAYER_S11_M10 `i_axi_AXI_W_LAYER_S11_M10
`endif 

`ifdef i_axi_AXI_W_LAYER_S11_M11
  `define AXI_W_LAYER_S11_M11 `i_axi_AXI_W_LAYER_S11_M11
`endif 

`ifdef i_axi_AXI_W_LAYER_S11_M12
  `define AXI_W_LAYER_S11_M12 `i_axi_AXI_W_LAYER_S11_M12
`endif 

`ifdef i_axi_AXI_W_LAYER_S11_M13
  `define AXI_W_LAYER_S11_M13 `i_axi_AXI_W_LAYER_S11_M13
`endif 

`ifdef i_axi_AXI_W_LAYER_S11_M14
  `define AXI_W_LAYER_S11_M14 `i_axi_AXI_W_LAYER_S11_M14
`endif 

`ifdef i_axi_AXI_W_LAYER_S11_M15
  `define AXI_W_LAYER_S11_M15 `i_axi_AXI_W_LAYER_S11_M15
`endif 

`ifdef i_axi_AXI_W_LAYER_S11_M16
  `define AXI_W_LAYER_S11_M16 `i_axi_AXI_W_LAYER_S11_M16
`endif 

`ifdef i_axi_AXI_AR_LAYER_S12_M1
  `define AXI_AR_LAYER_S12_M1 `i_axi_AXI_AR_LAYER_S12_M1
`endif 

`ifdef i_axi_AXI_AR_LAYER_S12_M2
  `define AXI_AR_LAYER_S12_M2 `i_axi_AXI_AR_LAYER_S12_M2
`endif 

`ifdef i_axi_AXI_AR_LAYER_S12_M3
  `define AXI_AR_LAYER_S12_M3 `i_axi_AXI_AR_LAYER_S12_M3
`endif 

`ifdef i_axi_AXI_AR_LAYER_S12_M4
  `define AXI_AR_LAYER_S12_M4 `i_axi_AXI_AR_LAYER_S12_M4
`endif 

`ifdef i_axi_AXI_AR_LAYER_S12_M5
  `define AXI_AR_LAYER_S12_M5 `i_axi_AXI_AR_LAYER_S12_M5
`endif 

`ifdef i_axi_AXI_AR_LAYER_S12_M6
  `define AXI_AR_LAYER_S12_M6 `i_axi_AXI_AR_LAYER_S12_M6
`endif 

`ifdef i_axi_AXI_AR_LAYER_S12_M7
  `define AXI_AR_LAYER_S12_M7 `i_axi_AXI_AR_LAYER_S12_M7
`endif 

`ifdef i_axi_AXI_AR_LAYER_S12_M8
  `define AXI_AR_LAYER_S12_M8 `i_axi_AXI_AR_LAYER_S12_M8
`endif 

`ifdef i_axi_AXI_AR_LAYER_S12_M9
  `define AXI_AR_LAYER_S12_M9 `i_axi_AXI_AR_LAYER_S12_M9
`endif 

`ifdef i_axi_AXI_AR_LAYER_S12_M10
  `define AXI_AR_LAYER_S12_M10 `i_axi_AXI_AR_LAYER_S12_M10
`endif 

`ifdef i_axi_AXI_AR_LAYER_S12_M11
  `define AXI_AR_LAYER_S12_M11 `i_axi_AXI_AR_LAYER_S12_M11
`endif 

`ifdef i_axi_AXI_AR_LAYER_S12_M12
  `define AXI_AR_LAYER_S12_M12 `i_axi_AXI_AR_LAYER_S12_M12
`endif 

`ifdef i_axi_AXI_AR_LAYER_S12_M13
  `define AXI_AR_LAYER_S12_M13 `i_axi_AXI_AR_LAYER_S12_M13
`endif 

`ifdef i_axi_AXI_AR_LAYER_S12_M14
  `define AXI_AR_LAYER_S12_M14 `i_axi_AXI_AR_LAYER_S12_M14
`endif 

`ifdef i_axi_AXI_AR_LAYER_S12_M15
  `define AXI_AR_LAYER_S12_M15 `i_axi_AXI_AR_LAYER_S12_M15
`endif 

`ifdef i_axi_AXI_AR_LAYER_S12_M16
  `define AXI_AR_LAYER_S12_M16 `i_axi_AXI_AR_LAYER_S12_M16
`endif 

`ifdef i_axi_AXI_AW_LAYER_S12_M1
  `define AXI_AW_LAYER_S12_M1 `i_axi_AXI_AW_LAYER_S12_M1
`endif 

`ifdef i_axi_AXI_AW_LAYER_S12_M2
  `define AXI_AW_LAYER_S12_M2 `i_axi_AXI_AW_LAYER_S12_M2
`endif 

`ifdef i_axi_AXI_AW_LAYER_S12_M3
  `define AXI_AW_LAYER_S12_M3 `i_axi_AXI_AW_LAYER_S12_M3
`endif 

`ifdef i_axi_AXI_AW_LAYER_S12_M4
  `define AXI_AW_LAYER_S12_M4 `i_axi_AXI_AW_LAYER_S12_M4
`endif 

`ifdef i_axi_AXI_AW_LAYER_S12_M5
  `define AXI_AW_LAYER_S12_M5 `i_axi_AXI_AW_LAYER_S12_M5
`endif 

`ifdef i_axi_AXI_AW_LAYER_S12_M6
  `define AXI_AW_LAYER_S12_M6 `i_axi_AXI_AW_LAYER_S12_M6
`endif 

`ifdef i_axi_AXI_AW_LAYER_S12_M7
  `define AXI_AW_LAYER_S12_M7 `i_axi_AXI_AW_LAYER_S12_M7
`endif 

`ifdef i_axi_AXI_AW_LAYER_S12_M8
  `define AXI_AW_LAYER_S12_M8 `i_axi_AXI_AW_LAYER_S12_M8
`endif 

`ifdef i_axi_AXI_AW_LAYER_S12_M9
  `define AXI_AW_LAYER_S12_M9 `i_axi_AXI_AW_LAYER_S12_M9
`endif 

`ifdef i_axi_AXI_AW_LAYER_S12_M10
  `define AXI_AW_LAYER_S12_M10 `i_axi_AXI_AW_LAYER_S12_M10
`endif 

`ifdef i_axi_AXI_AW_LAYER_S12_M11
  `define AXI_AW_LAYER_S12_M11 `i_axi_AXI_AW_LAYER_S12_M11
`endif 

`ifdef i_axi_AXI_AW_LAYER_S12_M12
  `define AXI_AW_LAYER_S12_M12 `i_axi_AXI_AW_LAYER_S12_M12
`endif 

`ifdef i_axi_AXI_AW_LAYER_S12_M13
  `define AXI_AW_LAYER_S12_M13 `i_axi_AXI_AW_LAYER_S12_M13
`endif 

`ifdef i_axi_AXI_AW_LAYER_S12_M14
  `define AXI_AW_LAYER_S12_M14 `i_axi_AXI_AW_LAYER_S12_M14
`endif 

`ifdef i_axi_AXI_AW_LAYER_S12_M15
  `define AXI_AW_LAYER_S12_M15 `i_axi_AXI_AW_LAYER_S12_M15
`endif 

`ifdef i_axi_AXI_AW_LAYER_S12_M16
  `define AXI_AW_LAYER_S12_M16 `i_axi_AXI_AW_LAYER_S12_M16
`endif 

`ifdef i_axi_AXI_W_LAYER_S12_M1
  `define AXI_W_LAYER_S12_M1 `i_axi_AXI_W_LAYER_S12_M1
`endif 

`ifdef i_axi_AXI_W_LAYER_S12_M2
  `define AXI_W_LAYER_S12_M2 `i_axi_AXI_W_LAYER_S12_M2
`endif 

`ifdef i_axi_AXI_W_LAYER_S12_M3
  `define AXI_W_LAYER_S12_M3 `i_axi_AXI_W_LAYER_S12_M3
`endif 

`ifdef i_axi_AXI_W_LAYER_S12_M4
  `define AXI_W_LAYER_S12_M4 `i_axi_AXI_W_LAYER_S12_M4
`endif 

`ifdef i_axi_AXI_W_LAYER_S12_M5
  `define AXI_W_LAYER_S12_M5 `i_axi_AXI_W_LAYER_S12_M5
`endif 

`ifdef i_axi_AXI_W_LAYER_S12_M6
  `define AXI_W_LAYER_S12_M6 `i_axi_AXI_W_LAYER_S12_M6
`endif 

`ifdef i_axi_AXI_W_LAYER_S12_M7
  `define AXI_W_LAYER_S12_M7 `i_axi_AXI_W_LAYER_S12_M7
`endif 

`ifdef i_axi_AXI_W_LAYER_S12_M8
  `define AXI_W_LAYER_S12_M8 `i_axi_AXI_W_LAYER_S12_M8
`endif 

`ifdef i_axi_AXI_W_LAYER_S12_M9
  `define AXI_W_LAYER_S12_M9 `i_axi_AXI_W_LAYER_S12_M9
`endif 

`ifdef i_axi_AXI_W_LAYER_S12_M10
  `define AXI_W_LAYER_S12_M10 `i_axi_AXI_W_LAYER_S12_M10
`endif 

`ifdef i_axi_AXI_W_LAYER_S12_M11
  `define AXI_W_LAYER_S12_M11 `i_axi_AXI_W_LAYER_S12_M11
`endif 

`ifdef i_axi_AXI_W_LAYER_S12_M12
  `define AXI_W_LAYER_S12_M12 `i_axi_AXI_W_LAYER_S12_M12
`endif 

`ifdef i_axi_AXI_W_LAYER_S12_M13
  `define AXI_W_LAYER_S12_M13 `i_axi_AXI_W_LAYER_S12_M13
`endif 

`ifdef i_axi_AXI_W_LAYER_S12_M14
  `define AXI_W_LAYER_S12_M14 `i_axi_AXI_W_LAYER_S12_M14
`endif 

`ifdef i_axi_AXI_W_LAYER_S12_M15
  `define AXI_W_LAYER_S12_M15 `i_axi_AXI_W_LAYER_S12_M15
`endif 

`ifdef i_axi_AXI_W_LAYER_S12_M16
  `define AXI_W_LAYER_S12_M16 `i_axi_AXI_W_LAYER_S12_M16
`endif 

`ifdef i_axi_AXI_AR_LAYER_S13_M1
  `define AXI_AR_LAYER_S13_M1 `i_axi_AXI_AR_LAYER_S13_M1
`endif 

`ifdef i_axi_AXI_AR_LAYER_S13_M2
  `define AXI_AR_LAYER_S13_M2 `i_axi_AXI_AR_LAYER_S13_M2
`endif 

`ifdef i_axi_AXI_AR_LAYER_S13_M3
  `define AXI_AR_LAYER_S13_M3 `i_axi_AXI_AR_LAYER_S13_M3
`endif 

`ifdef i_axi_AXI_AR_LAYER_S13_M4
  `define AXI_AR_LAYER_S13_M4 `i_axi_AXI_AR_LAYER_S13_M4
`endif 

`ifdef i_axi_AXI_AR_LAYER_S13_M5
  `define AXI_AR_LAYER_S13_M5 `i_axi_AXI_AR_LAYER_S13_M5
`endif 

`ifdef i_axi_AXI_AR_LAYER_S13_M6
  `define AXI_AR_LAYER_S13_M6 `i_axi_AXI_AR_LAYER_S13_M6
`endif 

`ifdef i_axi_AXI_AR_LAYER_S13_M7
  `define AXI_AR_LAYER_S13_M7 `i_axi_AXI_AR_LAYER_S13_M7
`endif 

`ifdef i_axi_AXI_AR_LAYER_S13_M8
  `define AXI_AR_LAYER_S13_M8 `i_axi_AXI_AR_LAYER_S13_M8
`endif 

`ifdef i_axi_AXI_AR_LAYER_S13_M9
  `define AXI_AR_LAYER_S13_M9 `i_axi_AXI_AR_LAYER_S13_M9
`endif 

`ifdef i_axi_AXI_AR_LAYER_S13_M10
  `define AXI_AR_LAYER_S13_M10 `i_axi_AXI_AR_LAYER_S13_M10
`endif 

`ifdef i_axi_AXI_AR_LAYER_S13_M11
  `define AXI_AR_LAYER_S13_M11 `i_axi_AXI_AR_LAYER_S13_M11
`endif 

`ifdef i_axi_AXI_AR_LAYER_S13_M12
  `define AXI_AR_LAYER_S13_M12 `i_axi_AXI_AR_LAYER_S13_M12
`endif 

`ifdef i_axi_AXI_AR_LAYER_S13_M13
  `define AXI_AR_LAYER_S13_M13 `i_axi_AXI_AR_LAYER_S13_M13
`endif 

`ifdef i_axi_AXI_AR_LAYER_S13_M14
  `define AXI_AR_LAYER_S13_M14 `i_axi_AXI_AR_LAYER_S13_M14
`endif 

`ifdef i_axi_AXI_AR_LAYER_S13_M15
  `define AXI_AR_LAYER_S13_M15 `i_axi_AXI_AR_LAYER_S13_M15
`endif 

`ifdef i_axi_AXI_AR_LAYER_S13_M16
  `define AXI_AR_LAYER_S13_M16 `i_axi_AXI_AR_LAYER_S13_M16
`endif 

`ifdef i_axi_AXI_AW_LAYER_S13_M1
  `define AXI_AW_LAYER_S13_M1 `i_axi_AXI_AW_LAYER_S13_M1
`endif 

`ifdef i_axi_AXI_AW_LAYER_S13_M2
  `define AXI_AW_LAYER_S13_M2 `i_axi_AXI_AW_LAYER_S13_M2
`endif 

`ifdef i_axi_AXI_AW_LAYER_S13_M3
  `define AXI_AW_LAYER_S13_M3 `i_axi_AXI_AW_LAYER_S13_M3
`endif 

`ifdef i_axi_AXI_AW_LAYER_S13_M4
  `define AXI_AW_LAYER_S13_M4 `i_axi_AXI_AW_LAYER_S13_M4
`endif 

`ifdef i_axi_AXI_AW_LAYER_S13_M5
  `define AXI_AW_LAYER_S13_M5 `i_axi_AXI_AW_LAYER_S13_M5
`endif 

`ifdef i_axi_AXI_AW_LAYER_S13_M6
  `define AXI_AW_LAYER_S13_M6 `i_axi_AXI_AW_LAYER_S13_M6
`endif 

`ifdef i_axi_AXI_AW_LAYER_S13_M7
  `define AXI_AW_LAYER_S13_M7 `i_axi_AXI_AW_LAYER_S13_M7
`endif 

`ifdef i_axi_AXI_AW_LAYER_S13_M8
  `define AXI_AW_LAYER_S13_M8 `i_axi_AXI_AW_LAYER_S13_M8
`endif 

`ifdef i_axi_AXI_AW_LAYER_S13_M9
  `define AXI_AW_LAYER_S13_M9 `i_axi_AXI_AW_LAYER_S13_M9
`endif 

`ifdef i_axi_AXI_AW_LAYER_S13_M10
  `define AXI_AW_LAYER_S13_M10 `i_axi_AXI_AW_LAYER_S13_M10
`endif 

`ifdef i_axi_AXI_AW_LAYER_S13_M11
  `define AXI_AW_LAYER_S13_M11 `i_axi_AXI_AW_LAYER_S13_M11
`endif 

`ifdef i_axi_AXI_AW_LAYER_S13_M12
  `define AXI_AW_LAYER_S13_M12 `i_axi_AXI_AW_LAYER_S13_M12
`endif 

`ifdef i_axi_AXI_AW_LAYER_S13_M13
  `define AXI_AW_LAYER_S13_M13 `i_axi_AXI_AW_LAYER_S13_M13
`endif 

`ifdef i_axi_AXI_AW_LAYER_S13_M14
  `define AXI_AW_LAYER_S13_M14 `i_axi_AXI_AW_LAYER_S13_M14
`endif 

`ifdef i_axi_AXI_AW_LAYER_S13_M15
  `define AXI_AW_LAYER_S13_M15 `i_axi_AXI_AW_LAYER_S13_M15
`endif 

`ifdef i_axi_AXI_AW_LAYER_S13_M16
  `define AXI_AW_LAYER_S13_M16 `i_axi_AXI_AW_LAYER_S13_M16
`endif 

`ifdef i_axi_AXI_W_LAYER_S13_M1
  `define AXI_W_LAYER_S13_M1 `i_axi_AXI_W_LAYER_S13_M1
`endif 

`ifdef i_axi_AXI_W_LAYER_S13_M2
  `define AXI_W_LAYER_S13_M2 `i_axi_AXI_W_LAYER_S13_M2
`endif 

`ifdef i_axi_AXI_W_LAYER_S13_M3
  `define AXI_W_LAYER_S13_M3 `i_axi_AXI_W_LAYER_S13_M3
`endif 

`ifdef i_axi_AXI_W_LAYER_S13_M4
  `define AXI_W_LAYER_S13_M4 `i_axi_AXI_W_LAYER_S13_M4
`endif 

`ifdef i_axi_AXI_W_LAYER_S13_M5
  `define AXI_W_LAYER_S13_M5 `i_axi_AXI_W_LAYER_S13_M5
`endif 

`ifdef i_axi_AXI_W_LAYER_S13_M6
  `define AXI_W_LAYER_S13_M6 `i_axi_AXI_W_LAYER_S13_M6
`endif 

`ifdef i_axi_AXI_W_LAYER_S13_M7
  `define AXI_W_LAYER_S13_M7 `i_axi_AXI_W_LAYER_S13_M7
`endif 

`ifdef i_axi_AXI_W_LAYER_S13_M8
  `define AXI_W_LAYER_S13_M8 `i_axi_AXI_W_LAYER_S13_M8
`endif 

`ifdef i_axi_AXI_W_LAYER_S13_M9
  `define AXI_W_LAYER_S13_M9 `i_axi_AXI_W_LAYER_S13_M9
`endif 

`ifdef i_axi_AXI_W_LAYER_S13_M10
  `define AXI_W_LAYER_S13_M10 `i_axi_AXI_W_LAYER_S13_M10
`endif 

`ifdef i_axi_AXI_W_LAYER_S13_M11
  `define AXI_W_LAYER_S13_M11 `i_axi_AXI_W_LAYER_S13_M11
`endif 

`ifdef i_axi_AXI_W_LAYER_S13_M12
  `define AXI_W_LAYER_S13_M12 `i_axi_AXI_W_LAYER_S13_M12
`endif 

`ifdef i_axi_AXI_W_LAYER_S13_M13
  `define AXI_W_LAYER_S13_M13 `i_axi_AXI_W_LAYER_S13_M13
`endif 

`ifdef i_axi_AXI_W_LAYER_S13_M14
  `define AXI_W_LAYER_S13_M14 `i_axi_AXI_W_LAYER_S13_M14
`endif 

`ifdef i_axi_AXI_W_LAYER_S13_M15
  `define AXI_W_LAYER_S13_M15 `i_axi_AXI_W_LAYER_S13_M15
`endif 

`ifdef i_axi_AXI_W_LAYER_S13_M16
  `define AXI_W_LAYER_S13_M16 `i_axi_AXI_W_LAYER_S13_M16
`endif 

`ifdef i_axi_AXI_AR_LAYER_S14_M1
  `define AXI_AR_LAYER_S14_M1 `i_axi_AXI_AR_LAYER_S14_M1
`endif 

`ifdef i_axi_AXI_AR_LAYER_S14_M2
  `define AXI_AR_LAYER_S14_M2 `i_axi_AXI_AR_LAYER_S14_M2
`endif 

`ifdef i_axi_AXI_AR_LAYER_S14_M3
  `define AXI_AR_LAYER_S14_M3 `i_axi_AXI_AR_LAYER_S14_M3
`endif 

`ifdef i_axi_AXI_AR_LAYER_S14_M4
  `define AXI_AR_LAYER_S14_M4 `i_axi_AXI_AR_LAYER_S14_M4
`endif 

`ifdef i_axi_AXI_AR_LAYER_S14_M5
  `define AXI_AR_LAYER_S14_M5 `i_axi_AXI_AR_LAYER_S14_M5
`endif 

`ifdef i_axi_AXI_AR_LAYER_S14_M6
  `define AXI_AR_LAYER_S14_M6 `i_axi_AXI_AR_LAYER_S14_M6
`endif 

`ifdef i_axi_AXI_AR_LAYER_S14_M7
  `define AXI_AR_LAYER_S14_M7 `i_axi_AXI_AR_LAYER_S14_M7
`endif 

`ifdef i_axi_AXI_AR_LAYER_S14_M8
  `define AXI_AR_LAYER_S14_M8 `i_axi_AXI_AR_LAYER_S14_M8
`endif 

`ifdef i_axi_AXI_AR_LAYER_S14_M9
  `define AXI_AR_LAYER_S14_M9 `i_axi_AXI_AR_LAYER_S14_M9
`endif 

`ifdef i_axi_AXI_AR_LAYER_S14_M10
  `define AXI_AR_LAYER_S14_M10 `i_axi_AXI_AR_LAYER_S14_M10
`endif 

`ifdef i_axi_AXI_AR_LAYER_S14_M11
  `define AXI_AR_LAYER_S14_M11 `i_axi_AXI_AR_LAYER_S14_M11
`endif 

`ifdef i_axi_AXI_AR_LAYER_S14_M12
  `define AXI_AR_LAYER_S14_M12 `i_axi_AXI_AR_LAYER_S14_M12
`endif 

`ifdef i_axi_AXI_AR_LAYER_S14_M13
  `define AXI_AR_LAYER_S14_M13 `i_axi_AXI_AR_LAYER_S14_M13
`endif 

`ifdef i_axi_AXI_AR_LAYER_S14_M14
  `define AXI_AR_LAYER_S14_M14 `i_axi_AXI_AR_LAYER_S14_M14
`endif 

`ifdef i_axi_AXI_AR_LAYER_S14_M15
  `define AXI_AR_LAYER_S14_M15 `i_axi_AXI_AR_LAYER_S14_M15
`endif 

`ifdef i_axi_AXI_AR_LAYER_S14_M16
  `define AXI_AR_LAYER_S14_M16 `i_axi_AXI_AR_LAYER_S14_M16
`endif 

`ifdef i_axi_AXI_AW_LAYER_S14_M1
  `define AXI_AW_LAYER_S14_M1 `i_axi_AXI_AW_LAYER_S14_M1
`endif 

`ifdef i_axi_AXI_AW_LAYER_S14_M2
  `define AXI_AW_LAYER_S14_M2 `i_axi_AXI_AW_LAYER_S14_M2
`endif 

`ifdef i_axi_AXI_AW_LAYER_S14_M3
  `define AXI_AW_LAYER_S14_M3 `i_axi_AXI_AW_LAYER_S14_M3
`endif 

`ifdef i_axi_AXI_AW_LAYER_S14_M4
  `define AXI_AW_LAYER_S14_M4 `i_axi_AXI_AW_LAYER_S14_M4
`endif 

`ifdef i_axi_AXI_AW_LAYER_S14_M5
  `define AXI_AW_LAYER_S14_M5 `i_axi_AXI_AW_LAYER_S14_M5
`endif 

`ifdef i_axi_AXI_AW_LAYER_S14_M6
  `define AXI_AW_LAYER_S14_M6 `i_axi_AXI_AW_LAYER_S14_M6
`endif 

`ifdef i_axi_AXI_AW_LAYER_S14_M7
  `define AXI_AW_LAYER_S14_M7 `i_axi_AXI_AW_LAYER_S14_M7
`endif 

`ifdef i_axi_AXI_AW_LAYER_S14_M8
  `define AXI_AW_LAYER_S14_M8 `i_axi_AXI_AW_LAYER_S14_M8
`endif 

`ifdef i_axi_AXI_AW_LAYER_S14_M9
  `define AXI_AW_LAYER_S14_M9 `i_axi_AXI_AW_LAYER_S14_M9
`endif 

`ifdef i_axi_AXI_AW_LAYER_S14_M10
  `define AXI_AW_LAYER_S14_M10 `i_axi_AXI_AW_LAYER_S14_M10
`endif 

`ifdef i_axi_AXI_AW_LAYER_S14_M11
  `define AXI_AW_LAYER_S14_M11 `i_axi_AXI_AW_LAYER_S14_M11
`endif 

`ifdef i_axi_AXI_AW_LAYER_S14_M12
  `define AXI_AW_LAYER_S14_M12 `i_axi_AXI_AW_LAYER_S14_M12
`endif 

`ifdef i_axi_AXI_AW_LAYER_S14_M13
  `define AXI_AW_LAYER_S14_M13 `i_axi_AXI_AW_LAYER_S14_M13
`endif 

`ifdef i_axi_AXI_AW_LAYER_S14_M14
  `define AXI_AW_LAYER_S14_M14 `i_axi_AXI_AW_LAYER_S14_M14
`endif 

`ifdef i_axi_AXI_AW_LAYER_S14_M15
  `define AXI_AW_LAYER_S14_M15 `i_axi_AXI_AW_LAYER_S14_M15
`endif 

`ifdef i_axi_AXI_AW_LAYER_S14_M16
  `define AXI_AW_LAYER_S14_M16 `i_axi_AXI_AW_LAYER_S14_M16
`endif 

`ifdef i_axi_AXI_W_LAYER_S14_M1
  `define AXI_W_LAYER_S14_M1 `i_axi_AXI_W_LAYER_S14_M1
`endif 

`ifdef i_axi_AXI_W_LAYER_S14_M2
  `define AXI_W_LAYER_S14_M2 `i_axi_AXI_W_LAYER_S14_M2
`endif 

`ifdef i_axi_AXI_W_LAYER_S14_M3
  `define AXI_W_LAYER_S14_M3 `i_axi_AXI_W_LAYER_S14_M3
`endif 

`ifdef i_axi_AXI_W_LAYER_S14_M4
  `define AXI_W_LAYER_S14_M4 `i_axi_AXI_W_LAYER_S14_M4
`endif 

`ifdef i_axi_AXI_W_LAYER_S14_M5
  `define AXI_W_LAYER_S14_M5 `i_axi_AXI_W_LAYER_S14_M5
`endif 

`ifdef i_axi_AXI_W_LAYER_S14_M6
  `define AXI_W_LAYER_S14_M6 `i_axi_AXI_W_LAYER_S14_M6
`endif 

`ifdef i_axi_AXI_W_LAYER_S14_M7
  `define AXI_W_LAYER_S14_M7 `i_axi_AXI_W_LAYER_S14_M7
`endif 

`ifdef i_axi_AXI_W_LAYER_S14_M8
  `define AXI_W_LAYER_S14_M8 `i_axi_AXI_W_LAYER_S14_M8
`endif 

`ifdef i_axi_AXI_W_LAYER_S14_M9
  `define AXI_W_LAYER_S14_M9 `i_axi_AXI_W_LAYER_S14_M9
`endif 

`ifdef i_axi_AXI_W_LAYER_S14_M10
  `define AXI_W_LAYER_S14_M10 `i_axi_AXI_W_LAYER_S14_M10
`endif 

`ifdef i_axi_AXI_W_LAYER_S14_M11
  `define AXI_W_LAYER_S14_M11 `i_axi_AXI_W_LAYER_S14_M11
`endif 

`ifdef i_axi_AXI_W_LAYER_S14_M12
  `define AXI_W_LAYER_S14_M12 `i_axi_AXI_W_LAYER_S14_M12
`endif 

`ifdef i_axi_AXI_W_LAYER_S14_M13
  `define AXI_W_LAYER_S14_M13 `i_axi_AXI_W_LAYER_S14_M13
`endif 

`ifdef i_axi_AXI_W_LAYER_S14_M14
  `define AXI_W_LAYER_S14_M14 `i_axi_AXI_W_LAYER_S14_M14
`endif 

`ifdef i_axi_AXI_W_LAYER_S14_M15
  `define AXI_W_LAYER_S14_M15 `i_axi_AXI_W_LAYER_S14_M15
`endif 

`ifdef i_axi_AXI_W_LAYER_S14_M16
  `define AXI_W_LAYER_S14_M16 `i_axi_AXI_W_LAYER_S14_M16
`endif 

`ifdef i_axi_AXI_AR_LAYER_S15_M1
  `define AXI_AR_LAYER_S15_M1 `i_axi_AXI_AR_LAYER_S15_M1
`endif 

`ifdef i_axi_AXI_AR_LAYER_S15_M2
  `define AXI_AR_LAYER_S15_M2 `i_axi_AXI_AR_LAYER_S15_M2
`endif 

`ifdef i_axi_AXI_AR_LAYER_S15_M3
  `define AXI_AR_LAYER_S15_M3 `i_axi_AXI_AR_LAYER_S15_M3
`endif 

`ifdef i_axi_AXI_AR_LAYER_S15_M4
  `define AXI_AR_LAYER_S15_M4 `i_axi_AXI_AR_LAYER_S15_M4
`endif 

`ifdef i_axi_AXI_AR_LAYER_S15_M5
  `define AXI_AR_LAYER_S15_M5 `i_axi_AXI_AR_LAYER_S15_M5
`endif 

`ifdef i_axi_AXI_AR_LAYER_S15_M6
  `define AXI_AR_LAYER_S15_M6 `i_axi_AXI_AR_LAYER_S15_M6
`endif 

`ifdef i_axi_AXI_AR_LAYER_S15_M7
  `define AXI_AR_LAYER_S15_M7 `i_axi_AXI_AR_LAYER_S15_M7
`endif 

`ifdef i_axi_AXI_AR_LAYER_S15_M8
  `define AXI_AR_LAYER_S15_M8 `i_axi_AXI_AR_LAYER_S15_M8
`endif 

`ifdef i_axi_AXI_AR_LAYER_S15_M9
  `define AXI_AR_LAYER_S15_M9 `i_axi_AXI_AR_LAYER_S15_M9
`endif 

`ifdef i_axi_AXI_AR_LAYER_S15_M10
  `define AXI_AR_LAYER_S15_M10 `i_axi_AXI_AR_LAYER_S15_M10
`endif 

`ifdef i_axi_AXI_AR_LAYER_S15_M11
  `define AXI_AR_LAYER_S15_M11 `i_axi_AXI_AR_LAYER_S15_M11
`endif 

`ifdef i_axi_AXI_AR_LAYER_S15_M12
  `define AXI_AR_LAYER_S15_M12 `i_axi_AXI_AR_LAYER_S15_M12
`endif 

`ifdef i_axi_AXI_AR_LAYER_S15_M13
  `define AXI_AR_LAYER_S15_M13 `i_axi_AXI_AR_LAYER_S15_M13
`endif 

`ifdef i_axi_AXI_AR_LAYER_S15_M14
  `define AXI_AR_LAYER_S15_M14 `i_axi_AXI_AR_LAYER_S15_M14
`endif 

`ifdef i_axi_AXI_AR_LAYER_S15_M15
  `define AXI_AR_LAYER_S15_M15 `i_axi_AXI_AR_LAYER_S15_M15
`endif 

`ifdef i_axi_AXI_AR_LAYER_S15_M16
  `define AXI_AR_LAYER_S15_M16 `i_axi_AXI_AR_LAYER_S15_M16
`endif 

`ifdef i_axi_AXI_AW_LAYER_S15_M1
  `define AXI_AW_LAYER_S15_M1 `i_axi_AXI_AW_LAYER_S15_M1
`endif 

`ifdef i_axi_AXI_AW_LAYER_S15_M2
  `define AXI_AW_LAYER_S15_M2 `i_axi_AXI_AW_LAYER_S15_M2
`endif 

`ifdef i_axi_AXI_AW_LAYER_S15_M3
  `define AXI_AW_LAYER_S15_M3 `i_axi_AXI_AW_LAYER_S15_M3
`endif 

`ifdef i_axi_AXI_AW_LAYER_S15_M4
  `define AXI_AW_LAYER_S15_M4 `i_axi_AXI_AW_LAYER_S15_M4
`endif 

`ifdef i_axi_AXI_AW_LAYER_S15_M5
  `define AXI_AW_LAYER_S15_M5 `i_axi_AXI_AW_LAYER_S15_M5
`endif 

`ifdef i_axi_AXI_AW_LAYER_S15_M6
  `define AXI_AW_LAYER_S15_M6 `i_axi_AXI_AW_LAYER_S15_M6
`endif 

`ifdef i_axi_AXI_AW_LAYER_S15_M7
  `define AXI_AW_LAYER_S15_M7 `i_axi_AXI_AW_LAYER_S15_M7
`endif 

`ifdef i_axi_AXI_AW_LAYER_S15_M8
  `define AXI_AW_LAYER_S15_M8 `i_axi_AXI_AW_LAYER_S15_M8
`endif 

`ifdef i_axi_AXI_AW_LAYER_S15_M9
  `define AXI_AW_LAYER_S15_M9 `i_axi_AXI_AW_LAYER_S15_M9
`endif 

`ifdef i_axi_AXI_AW_LAYER_S15_M10
  `define AXI_AW_LAYER_S15_M10 `i_axi_AXI_AW_LAYER_S15_M10
`endif 

`ifdef i_axi_AXI_AW_LAYER_S15_M11
  `define AXI_AW_LAYER_S15_M11 `i_axi_AXI_AW_LAYER_S15_M11
`endif 

`ifdef i_axi_AXI_AW_LAYER_S15_M12
  `define AXI_AW_LAYER_S15_M12 `i_axi_AXI_AW_LAYER_S15_M12
`endif 

`ifdef i_axi_AXI_AW_LAYER_S15_M13
  `define AXI_AW_LAYER_S15_M13 `i_axi_AXI_AW_LAYER_S15_M13
`endif 

`ifdef i_axi_AXI_AW_LAYER_S15_M14
  `define AXI_AW_LAYER_S15_M14 `i_axi_AXI_AW_LAYER_S15_M14
`endif 

`ifdef i_axi_AXI_AW_LAYER_S15_M15
  `define AXI_AW_LAYER_S15_M15 `i_axi_AXI_AW_LAYER_S15_M15
`endif 

`ifdef i_axi_AXI_AW_LAYER_S15_M16
  `define AXI_AW_LAYER_S15_M16 `i_axi_AXI_AW_LAYER_S15_M16
`endif 

`ifdef i_axi_AXI_W_LAYER_S15_M1
  `define AXI_W_LAYER_S15_M1 `i_axi_AXI_W_LAYER_S15_M1
`endif 

`ifdef i_axi_AXI_W_LAYER_S15_M2
  `define AXI_W_LAYER_S15_M2 `i_axi_AXI_W_LAYER_S15_M2
`endif 

`ifdef i_axi_AXI_W_LAYER_S15_M3
  `define AXI_W_LAYER_S15_M3 `i_axi_AXI_W_LAYER_S15_M3
`endif 

`ifdef i_axi_AXI_W_LAYER_S15_M4
  `define AXI_W_LAYER_S15_M4 `i_axi_AXI_W_LAYER_S15_M4
`endif 

`ifdef i_axi_AXI_W_LAYER_S15_M5
  `define AXI_W_LAYER_S15_M5 `i_axi_AXI_W_LAYER_S15_M5
`endif 

`ifdef i_axi_AXI_W_LAYER_S15_M6
  `define AXI_W_LAYER_S15_M6 `i_axi_AXI_W_LAYER_S15_M6
`endif 

`ifdef i_axi_AXI_W_LAYER_S15_M7
  `define AXI_W_LAYER_S15_M7 `i_axi_AXI_W_LAYER_S15_M7
`endif 

`ifdef i_axi_AXI_W_LAYER_S15_M8
  `define AXI_W_LAYER_S15_M8 `i_axi_AXI_W_LAYER_S15_M8
`endif 

`ifdef i_axi_AXI_W_LAYER_S15_M9
  `define AXI_W_LAYER_S15_M9 `i_axi_AXI_W_LAYER_S15_M9
`endif 

`ifdef i_axi_AXI_W_LAYER_S15_M10
  `define AXI_W_LAYER_S15_M10 `i_axi_AXI_W_LAYER_S15_M10
`endif 

`ifdef i_axi_AXI_W_LAYER_S15_M11
  `define AXI_W_LAYER_S15_M11 `i_axi_AXI_W_LAYER_S15_M11
`endif 

`ifdef i_axi_AXI_W_LAYER_S15_M12
  `define AXI_W_LAYER_S15_M12 `i_axi_AXI_W_LAYER_S15_M12
`endif 

`ifdef i_axi_AXI_W_LAYER_S15_M13
  `define AXI_W_LAYER_S15_M13 `i_axi_AXI_W_LAYER_S15_M13
`endif 

`ifdef i_axi_AXI_W_LAYER_S15_M14
  `define AXI_W_LAYER_S15_M14 `i_axi_AXI_W_LAYER_S15_M14
`endif 

`ifdef i_axi_AXI_W_LAYER_S15_M15
  `define AXI_W_LAYER_S15_M15 `i_axi_AXI_W_LAYER_S15_M15
`endif 

`ifdef i_axi_AXI_W_LAYER_S15_M16
  `define AXI_W_LAYER_S15_M16 `i_axi_AXI_W_LAYER_S15_M16
`endif 

`ifdef i_axi_AXI_AR_LAYER_S16_M1
  `define AXI_AR_LAYER_S16_M1 `i_axi_AXI_AR_LAYER_S16_M1
`endif 

`ifdef i_axi_AXI_AR_LAYER_S16_M2
  `define AXI_AR_LAYER_S16_M2 `i_axi_AXI_AR_LAYER_S16_M2
`endif 

`ifdef i_axi_AXI_AR_LAYER_S16_M3
  `define AXI_AR_LAYER_S16_M3 `i_axi_AXI_AR_LAYER_S16_M3
`endif 

`ifdef i_axi_AXI_AR_LAYER_S16_M4
  `define AXI_AR_LAYER_S16_M4 `i_axi_AXI_AR_LAYER_S16_M4
`endif 

`ifdef i_axi_AXI_AR_LAYER_S16_M5
  `define AXI_AR_LAYER_S16_M5 `i_axi_AXI_AR_LAYER_S16_M5
`endif 

`ifdef i_axi_AXI_AR_LAYER_S16_M6
  `define AXI_AR_LAYER_S16_M6 `i_axi_AXI_AR_LAYER_S16_M6
`endif 

`ifdef i_axi_AXI_AR_LAYER_S16_M7
  `define AXI_AR_LAYER_S16_M7 `i_axi_AXI_AR_LAYER_S16_M7
`endif 

`ifdef i_axi_AXI_AR_LAYER_S16_M8
  `define AXI_AR_LAYER_S16_M8 `i_axi_AXI_AR_LAYER_S16_M8
`endif 

`ifdef i_axi_AXI_AR_LAYER_S16_M9
  `define AXI_AR_LAYER_S16_M9 `i_axi_AXI_AR_LAYER_S16_M9
`endif 

`ifdef i_axi_AXI_AR_LAYER_S16_M10
  `define AXI_AR_LAYER_S16_M10 `i_axi_AXI_AR_LAYER_S16_M10
`endif 

`ifdef i_axi_AXI_AR_LAYER_S16_M11
  `define AXI_AR_LAYER_S16_M11 `i_axi_AXI_AR_LAYER_S16_M11
`endif 

`ifdef i_axi_AXI_AR_LAYER_S16_M12
  `define AXI_AR_LAYER_S16_M12 `i_axi_AXI_AR_LAYER_S16_M12
`endif 

`ifdef i_axi_AXI_AR_LAYER_S16_M13
  `define AXI_AR_LAYER_S16_M13 `i_axi_AXI_AR_LAYER_S16_M13
`endif 

`ifdef i_axi_AXI_AR_LAYER_S16_M14
  `define AXI_AR_LAYER_S16_M14 `i_axi_AXI_AR_LAYER_S16_M14
`endif 

`ifdef i_axi_AXI_AR_LAYER_S16_M15
  `define AXI_AR_LAYER_S16_M15 `i_axi_AXI_AR_LAYER_S16_M15
`endif 

`ifdef i_axi_AXI_AR_LAYER_S16_M16
  `define AXI_AR_LAYER_S16_M16 `i_axi_AXI_AR_LAYER_S16_M16
`endif 

`ifdef i_axi_AXI_AW_LAYER_S16_M1
  `define AXI_AW_LAYER_S16_M1 `i_axi_AXI_AW_LAYER_S16_M1
`endif 

`ifdef i_axi_AXI_AW_LAYER_S16_M2
  `define AXI_AW_LAYER_S16_M2 `i_axi_AXI_AW_LAYER_S16_M2
`endif 

`ifdef i_axi_AXI_AW_LAYER_S16_M3
  `define AXI_AW_LAYER_S16_M3 `i_axi_AXI_AW_LAYER_S16_M3
`endif 

`ifdef i_axi_AXI_AW_LAYER_S16_M4
  `define AXI_AW_LAYER_S16_M4 `i_axi_AXI_AW_LAYER_S16_M4
`endif 

`ifdef i_axi_AXI_AW_LAYER_S16_M5
  `define AXI_AW_LAYER_S16_M5 `i_axi_AXI_AW_LAYER_S16_M5
`endif 

`ifdef i_axi_AXI_AW_LAYER_S16_M6
  `define AXI_AW_LAYER_S16_M6 `i_axi_AXI_AW_LAYER_S16_M6
`endif 

`ifdef i_axi_AXI_AW_LAYER_S16_M7
  `define AXI_AW_LAYER_S16_M7 `i_axi_AXI_AW_LAYER_S16_M7
`endif 

`ifdef i_axi_AXI_AW_LAYER_S16_M8
  `define AXI_AW_LAYER_S16_M8 `i_axi_AXI_AW_LAYER_S16_M8
`endif 

`ifdef i_axi_AXI_AW_LAYER_S16_M9
  `define AXI_AW_LAYER_S16_M9 `i_axi_AXI_AW_LAYER_S16_M9
`endif 

`ifdef i_axi_AXI_AW_LAYER_S16_M10
  `define AXI_AW_LAYER_S16_M10 `i_axi_AXI_AW_LAYER_S16_M10
`endif 

`ifdef i_axi_AXI_AW_LAYER_S16_M11
  `define AXI_AW_LAYER_S16_M11 `i_axi_AXI_AW_LAYER_S16_M11
`endif 

`ifdef i_axi_AXI_AW_LAYER_S16_M12
  `define AXI_AW_LAYER_S16_M12 `i_axi_AXI_AW_LAYER_S16_M12
`endif 

`ifdef i_axi_AXI_AW_LAYER_S16_M13
  `define AXI_AW_LAYER_S16_M13 `i_axi_AXI_AW_LAYER_S16_M13
`endif 

`ifdef i_axi_AXI_AW_LAYER_S16_M14
  `define AXI_AW_LAYER_S16_M14 `i_axi_AXI_AW_LAYER_S16_M14
`endif 

`ifdef i_axi_AXI_AW_LAYER_S16_M15
  `define AXI_AW_LAYER_S16_M15 `i_axi_AXI_AW_LAYER_S16_M15
`endif 

`ifdef i_axi_AXI_AW_LAYER_S16_M16
  `define AXI_AW_LAYER_S16_M16 `i_axi_AXI_AW_LAYER_S16_M16
`endif 

`ifdef i_axi_AXI_W_LAYER_S16_M1
  `define AXI_W_LAYER_S16_M1 `i_axi_AXI_W_LAYER_S16_M1
`endif 

`ifdef i_axi_AXI_W_LAYER_S16_M2
  `define AXI_W_LAYER_S16_M2 `i_axi_AXI_W_LAYER_S16_M2
`endif 

`ifdef i_axi_AXI_W_LAYER_S16_M3
  `define AXI_W_LAYER_S16_M3 `i_axi_AXI_W_LAYER_S16_M3
`endif 

`ifdef i_axi_AXI_W_LAYER_S16_M4
  `define AXI_W_LAYER_S16_M4 `i_axi_AXI_W_LAYER_S16_M4
`endif 

`ifdef i_axi_AXI_W_LAYER_S16_M5
  `define AXI_W_LAYER_S16_M5 `i_axi_AXI_W_LAYER_S16_M5
`endif 

`ifdef i_axi_AXI_W_LAYER_S16_M6
  `define AXI_W_LAYER_S16_M6 `i_axi_AXI_W_LAYER_S16_M6
`endif 

`ifdef i_axi_AXI_W_LAYER_S16_M7
  `define AXI_W_LAYER_S16_M7 `i_axi_AXI_W_LAYER_S16_M7
`endif 

`ifdef i_axi_AXI_W_LAYER_S16_M8
  `define AXI_W_LAYER_S16_M8 `i_axi_AXI_W_LAYER_S16_M8
`endif 

`ifdef i_axi_AXI_W_LAYER_S16_M9
  `define AXI_W_LAYER_S16_M9 `i_axi_AXI_W_LAYER_S16_M9
`endif 

`ifdef i_axi_AXI_W_LAYER_S16_M10
  `define AXI_W_LAYER_S16_M10 `i_axi_AXI_W_LAYER_S16_M10
`endif 

`ifdef i_axi_AXI_W_LAYER_S16_M11
  `define AXI_W_LAYER_S16_M11 `i_axi_AXI_W_LAYER_S16_M11
`endif 

`ifdef i_axi_AXI_W_LAYER_S16_M12
  `define AXI_W_LAYER_S16_M12 `i_axi_AXI_W_LAYER_S16_M12
`endif 

`ifdef i_axi_AXI_W_LAYER_S16_M13
  `define AXI_W_LAYER_S16_M13 `i_axi_AXI_W_LAYER_S16_M13
`endif 

`ifdef i_axi_AXI_W_LAYER_S16_M14
  `define AXI_W_LAYER_S16_M14 `i_axi_AXI_W_LAYER_S16_M14
`endif 

`ifdef i_axi_AXI_W_LAYER_S16_M15
  `define AXI_W_LAYER_S16_M15 `i_axi_AXI_W_LAYER_S16_M15
`endif 

`ifdef i_axi_AXI_W_LAYER_S16_M16
  `define AXI_W_LAYER_S16_M16 `i_axi_AXI_W_LAYER_S16_M16
`endif 

`ifdef i_axi_AXI_ALL_R_LAYER_SHARED
  `define AXI_ALL_R_LAYER_SHARED `i_axi_AXI_ALL_R_LAYER_SHARED
`endif 

`ifdef i_axi_AXI_R_LAYER_M1_S0
  `define AXI_R_LAYER_M1_S0 `i_axi_AXI_R_LAYER_M1_S0
`endif 

`ifdef i_axi_AXI_R_LAYER_M1_S1
  `define AXI_R_LAYER_M1_S1 `i_axi_AXI_R_LAYER_M1_S1
`endif 

`ifdef i_axi_AXI_R_LAYER_M1_S2
  `define AXI_R_LAYER_M1_S2 `i_axi_AXI_R_LAYER_M1_S2
`endif 

`ifdef i_axi_AXI_R_LAYER_M1_S3
  `define AXI_R_LAYER_M1_S3 `i_axi_AXI_R_LAYER_M1_S3
`endif 

`ifdef i_axi_AXI_R_LAYER_M1_S4
  `define AXI_R_LAYER_M1_S4 `i_axi_AXI_R_LAYER_M1_S4
`endif 

`ifdef i_axi_AXI_R_LAYER_M1_S5
  `define AXI_R_LAYER_M1_S5 `i_axi_AXI_R_LAYER_M1_S5
`endif 

`ifdef i_axi_AXI_R_LAYER_M1_S6
  `define AXI_R_LAYER_M1_S6 `i_axi_AXI_R_LAYER_M1_S6
`endif 

`ifdef i_axi_AXI_R_LAYER_M1_S7
  `define AXI_R_LAYER_M1_S7 `i_axi_AXI_R_LAYER_M1_S7
`endif 

`ifdef i_axi_AXI_R_LAYER_M1_S8
  `define AXI_R_LAYER_M1_S8 `i_axi_AXI_R_LAYER_M1_S8
`endif 

`ifdef i_axi_AXI_R_LAYER_M1_S9
  `define AXI_R_LAYER_M1_S9 `i_axi_AXI_R_LAYER_M1_S9
`endif 

`ifdef i_axi_AXI_R_LAYER_M1_S10
  `define AXI_R_LAYER_M1_S10 `i_axi_AXI_R_LAYER_M1_S10
`endif 

`ifdef i_axi_AXI_R_LAYER_M1_S11
  `define AXI_R_LAYER_M1_S11 `i_axi_AXI_R_LAYER_M1_S11
`endif 

`ifdef i_axi_AXI_R_LAYER_M1_S12
  `define AXI_R_LAYER_M1_S12 `i_axi_AXI_R_LAYER_M1_S12
`endif 

`ifdef i_axi_AXI_R_LAYER_M1_S13
  `define AXI_R_LAYER_M1_S13 `i_axi_AXI_R_LAYER_M1_S13
`endif 

`ifdef i_axi_AXI_R_LAYER_M1_S14
  `define AXI_R_LAYER_M1_S14 `i_axi_AXI_R_LAYER_M1_S14
`endif 

`ifdef i_axi_AXI_R_LAYER_M1_S15
  `define AXI_R_LAYER_M1_S15 `i_axi_AXI_R_LAYER_M1_S15
`endif 

`ifdef i_axi_AXI_R_LAYER_M1_S16
  `define AXI_R_LAYER_M1_S16 `i_axi_AXI_R_LAYER_M1_S16
`endif 

`ifdef i_axi_AXI_ALL_B_LAYER_SHARED
  `define AXI_ALL_B_LAYER_SHARED `i_axi_AXI_ALL_B_LAYER_SHARED
`endif 

`ifdef i_axi_AXI_B_LAYER_M1_S0
  `define AXI_B_LAYER_M1_S0 `i_axi_AXI_B_LAYER_M1_S0
`endif 

`ifdef i_axi_AXI_B_LAYER_M1_S1
  `define AXI_B_LAYER_M1_S1 `i_axi_AXI_B_LAYER_M1_S1
`endif 

`ifdef i_axi_AXI_B_LAYER_M1_S2
  `define AXI_B_LAYER_M1_S2 `i_axi_AXI_B_LAYER_M1_S2
`endif 

`ifdef i_axi_AXI_B_LAYER_M1_S3
  `define AXI_B_LAYER_M1_S3 `i_axi_AXI_B_LAYER_M1_S3
`endif 

`ifdef i_axi_AXI_B_LAYER_M1_S4
  `define AXI_B_LAYER_M1_S4 `i_axi_AXI_B_LAYER_M1_S4
`endif 

`ifdef i_axi_AXI_B_LAYER_M1_S5
  `define AXI_B_LAYER_M1_S5 `i_axi_AXI_B_LAYER_M1_S5
`endif 

`ifdef i_axi_AXI_B_LAYER_M1_S6
  `define AXI_B_LAYER_M1_S6 `i_axi_AXI_B_LAYER_M1_S6
`endif 

`ifdef i_axi_AXI_B_LAYER_M1_S7
  `define AXI_B_LAYER_M1_S7 `i_axi_AXI_B_LAYER_M1_S7
`endif 

`ifdef i_axi_AXI_B_LAYER_M1_S8
  `define AXI_B_LAYER_M1_S8 `i_axi_AXI_B_LAYER_M1_S8
`endif 

`ifdef i_axi_AXI_B_LAYER_M1_S9
  `define AXI_B_LAYER_M1_S9 `i_axi_AXI_B_LAYER_M1_S9
`endif 

`ifdef i_axi_AXI_B_LAYER_M1_S10
  `define AXI_B_LAYER_M1_S10 `i_axi_AXI_B_LAYER_M1_S10
`endif 

`ifdef i_axi_AXI_B_LAYER_M1_S11
  `define AXI_B_LAYER_M1_S11 `i_axi_AXI_B_LAYER_M1_S11
`endif 

`ifdef i_axi_AXI_B_LAYER_M1_S12
  `define AXI_B_LAYER_M1_S12 `i_axi_AXI_B_LAYER_M1_S12
`endif 

`ifdef i_axi_AXI_B_LAYER_M1_S13
  `define AXI_B_LAYER_M1_S13 `i_axi_AXI_B_LAYER_M1_S13
`endif 

`ifdef i_axi_AXI_B_LAYER_M1_S14
  `define AXI_B_LAYER_M1_S14 `i_axi_AXI_B_LAYER_M1_S14
`endif 

`ifdef i_axi_AXI_B_LAYER_M1_S15
  `define AXI_B_LAYER_M1_S15 `i_axi_AXI_B_LAYER_M1_S15
`endif 

`ifdef i_axi_AXI_B_LAYER_M1_S16
  `define AXI_B_LAYER_M1_S16 `i_axi_AXI_B_LAYER_M1_S16
`endif 

`ifdef i_axi_AXI_R_LAYER_M2_S0
  `define AXI_R_LAYER_M2_S0 `i_axi_AXI_R_LAYER_M2_S0
`endif 

`ifdef i_axi_AXI_R_LAYER_M2_S1
  `define AXI_R_LAYER_M2_S1 `i_axi_AXI_R_LAYER_M2_S1
`endif 

`ifdef i_axi_AXI_R_LAYER_M2_S2
  `define AXI_R_LAYER_M2_S2 `i_axi_AXI_R_LAYER_M2_S2
`endif 

`ifdef i_axi_AXI_R_LAYER_M2_S3
  `define AXI_R_LAYER_M2_S3 `i_axi_AXI_R_LAYER_M2_S3
`endif 

`ifdef i_axi_AXI_R_LAYER_M2_S4
  `define AXI_R_LAYER_M2_S4 `i_axi_AXI_R_LAYER_M2_S4
`endif 

`ifdef i_axi_AXI_R_LAYER_M2_S5
  `define AXI_R_LAYER_M2_S5 `i_axi_AXI_R_LAYER_M2_S5
`endif 

`ifdef i_axi_AXI_R_LAYER_M2_S6
  `define AXI_R_LAYER_M2_S6 `i_axi_AXI_R_LAYER_M2_S6
`endif 

`ifdef i_axi_AXI_R_LAYER_M2_S7
  `define AXI_R_LAYER_M2_S7 `i_axi_AXI_R_LAYER_M2_S7
`endif 

`ifdef i_axi_AXI_R_LAYER_M2_S8
  `define AXI_R_LAYER_M2_S8 `i_axi_AXI_R_LAYER_M2_S8
`endif 

`ifdef i_axi_AXI_R_LAYER_M2_S9
  `define AXI_R_LAYER_M2_S9 `i_axi_AXI_R_LAYER_M2_S9
`endif 

`ifdef i_axi_AXI_R_LAYER_M2_S10
  `define AXI_R_LAYER_M2_S10 `i_axi_AXI_R_LAYER_M2_S10
`endif 

`ifdef i_axi_AXI_R_LAYER_M2_S11
  `define AXI_R_LAYER_M2_S11 `i_axi_AXI_R_LAYER_M2_S11
`endif 

`ifdef i_axi_AXI_R_LAYER_M2_S12
  `define AXI_R_LAYER_M2_S12 `i_axi_AXI_R_LAYER_M2_S12
`endif 

`ifdef i_axi_AXI_R_LAYER_M2_S13
  `define AXI_R_LAYER_M2_S13 `i_axi_AXI_R_LAYER_M2_S13
`endif 

`ifdef i_axi_AXI_R_LAYER_M2_S14
  `define AXI_R_LAYER_M2_S14 `i_axi_AXI_R_LAYER_M2_S14
`endif 

`ifdef i_axi_AXI_R_LAYER_M2_S15
  `define AXI_R_LAYER_M2_S15 `i_axi_AXI_R_LAYER_M2_S15
`endif 

`ifdef i_axi_AXI_R_LAYER_M2_S16
  `define AXI_R_LAYER_M2_S16 `i_axi_AXI_R_LAYER_M2_S16
`endif 

`ifdef i_axi_AXI_B_LAYER_M2_S0
  `define AXI_B_LAYER_M2_S0 `i_axi_AXI_B_LAYER_M2_S0
`endif 

`ifdef i_axi_AXI_B_LAYER_M2_S1
  `define AXI_B_LAYER_M2_S1 `i_axi_AXI_B_LAYER_M2_S1
`endif 

`ifdef i_axi_AXI_B_LAYER_M2_S2
  `define AXI_B_LAYER_M2_S2 `i_axi_AXI_B_LAYER_M2_S2
`endif 

`ifdef i_axi_AXI_B_LAYER_M2_S3
  `define AXI_B_LAYER_M2_S3 `i_axi_AXI_B_LAYER_M2_S3
`endif 

`ifdef i_axi_AXI_B_LAYER_M2_S4
  `define AXI_B_LAYER_M2_S4 `i_axi_AXI_B_LAYER_M2_S4
`endif 

`ifdef i_axi_AXI_B_LAYER_M2_S5
  `define AXI_B_LAYER_M2_S5 `i_axi_AXI_B_LAYER_M2_S5
`endif 

`ifdef i_axi_AXI_B_LAYER_M2_S6
  `define AXI_B_LAYER_M2_S6 `i_axi_AXI_B_LAYER_M2_S6
`endif 

`ifdef i_axi_AXI_B_LAYER_M2_S7
  `define AXI_B_LAYER_M2_S7 `i_axi_AXI_B_LAYER_M2_S7
`endif 

`ifdef i_axi_AXI_B_LAYER_M2_S8
  `define AXI_B_LAYER_M2_S8 `i_axi_AXI_B_LAYER_M2_S8
`endif 

`ifdef i_axi_AXI_B_LAYER_M2_S9
  `define AXI_B_LAYER_M2_S9 `i_axi_AXI_B_LAYER_M2_S9
`endif 

`ifdef i_axi_AXI_B_LAYER_M2_S10
  `define AXI_B_LAYER_M2_S10 `i_axi_AXI_B_LAYER_M2_S10
`endif 

`ifdef i_axi_AXI_B_LAYER_M2_S11
  `define AXI_B_LAYER_M2_S11 `i_axi_AXI_B_LAYER_M2_S11
`endif 

`ifdef i_axi_AXI_B_LAYER_M2_S12
  `define AXI_B_LAYER_M2_S12 `i_axi_AXI_B_LAYER_M2_S12
`endif 

`ifdef i_axi_AXI_B_LAYER_M2_S13
  `define AXI_B_LAYER_M2_S13 `i_axi_AXI_B_LAYER_M2_S13
`endif 

`ifdef i_axi_AXI_B_LAYER_M2_S14
  `define AXI_B_LAYER_M2_S14 `i_axi_AXI_B_LAYER_M2_S14
`endif 

`ifdef i_axi_AXI_B_LAYER_M2_S15
  `define AXI_B_LAYER_M2_S15 `i_axi_AXI_B_LAYER_M2_S15
`endif 

`ifdef i_axi_AXI_B_LAYER_M2_S16
  `define AXI_B_LAYER_M2_S16 `i_axi_AXI_B_LAYER_M2_S16
`endif 

`ifdef i_axi_AXI_R_LAYER_M3_S0
  `define AXI_R_LAYER_M3_S0 `i_axi_AXI_R_LAYER_M3_S0
`endif 

`ifdef i_axi_AXI_R_LAYER_M3_S1
  `define AXI_R_LAYER_M3_S1 `i_axi_AXI_R_LAYER_M3_S1
`endif 

`ifdef i_axi_AXI_R_LAYER_M3_S2
  `define AXI_R_LAYER_M3_S2 `i_axi_AXI_R_LAYER_M3_S2
`endif 

`ifdef i_axi_AXI_R_LAYER_M3_S3
  `define AXI_R_LAYER_M3_S3 `i_axi_AXI_R_LAYER_M3_S3
`endif 

`ifdef i_axi_AXI_R_LAYER_M3_S4
  `define AXI_R_LAYER_M3_S4 `i_axi_AXI_R_LAYER_M3_S4
`endif 

`ifdef i_axi_AXI_R_LAYER_M3_S5
  `define AXI_R_LAYER_M3_S5 `i_axi_AXI_R_LAYER_M3_S5
`endif 

`ifdef i_axi_AXI_R_LAYER_M3_S6
  `define AXI_R_LAYER_M3_S6 `i_axi_AXI_R_LAYER_M3_S6
`endif 

`ifdef i_axi_AXI_R_LAYER_M3_S7
  `define AXI_R_LAYER_M3_S7 `i_axi_AXI_R_LAYER_M3_S7
`endif 

`ifdef i_axi_AXI_R_LAYER_M3_S8
  `define AXI_R_LAYER_M3_S8 `i_axi_AXI_R_LAYER_M3_S8
`endif 

`ifdef i_axi_AXI_R_LAYER_M3_S9
  `define AXI_R_LAYER_M3_S9 `i_axi_AXI_R_LAYER_M3_S9
`endif 

`ifdef i_axi_AXI_R_LAYER_M3_S10
  `define AXI_R_LAYER_M3_S10 `i_axi_AXI_R_LAYER_M3_S10
`endif 

`ifdef i_axi_AXI_R_LAYER_M3_S11
  `define AXI_R_LAYER_M3_S11 `i_axi_AXI_R_LAYER_M3_S11
`endif 

`ifdef i_axi_AXI_R_LAYER_M3_S12
  `define AXI_R_LAYER_M3_S12 `i_axi_AXI_R_LAYER_M3_S12
`endif 

`ifdef i_axi_AXI_R_LAYER_M3_S13
  `define AXI_R_LAYER_M3_S13 `i_axi_AXI_R_LAYER_M3_S13
`endif 

`ifdef i_axi_AXI_R_LAYER_M3_S14
  `define AXI_R_LAYER_M3_S14 `i_axi_AXI_R_LAYER_M3_S14
`endif 

`ifdef i_axi_AXI_R_LAYER_M3_S15
  `define AXI_R_LAYER_M3_S15 `i_axi_AXI_R_LAYER_M3_S15
`endif 

`ifdef i_axi_AXI_R_LAYER_M3_S16
  `define AXI_R_LAYER_M3_S16 `i_axi_AXI_R_LAYER_M3_S16
`endif 

`ifdef i_axi_AXI_B_LAYER_M3_S0
  `define AXI_B_LAYER_M3_S0 `i_axi_AXI_B_LAYER_M3_S0
`endif 

`ifdef i_axi_AXI_B_LAYER_M3_S1
  `define AXI_B_LAYER_M3_S1 `i_axi_AXI_B_LAYER_M3_S1
`endif 

`ifdef i_axi_AXI_B_LAYER_M3_S2
  `define AXI_B_LAYER_M3_S2 `i_axi_AXI_B_LAYER_M3_S2
`endif 

`ifdef i_axi_AXI_B_LAYER_M3_S3
  `define AXI_B_LAYER_M3_S3 `i_axi_AXI_B_LAYER_M3_S3
`endif 

`ifdef i_axi_AXI_B_LAYER_M3_S4
  `define AXI_B_LAYER_M3_S4 `i_axi_AXI_B_LAYER_M3_S4
`endif 

`ifdef i_axi_AXI_B_LAYER_M3_S5
  `define AXI_B_LAYER_M3_S5 `i_axi_AXI_B_LAYER_M3_S5
`endif 

`ifdef i_axi_AXI_B_LAYER_M3_S6
  `define AXI_B_LAYER_M3_S6 `i_axi_AXI_B_LAYER_M3_S6
`endif 

`ifdef i_axi_AXI_B_LAYER_M3_S7
  `define AXI_B_LAYER_M3_S7 `i_axi_AXI_B_LAYER_M3_S7
`endif 

`ifdef i_axi_AXI_B_LAYER_M3_S8
  `define AXI_B_LAYER_M3_S8 `i_axi_AXI_B_LAYER_M3_S8
`endif 

`ifdef i_axi_AXI_B_LAYER_M3_S9
  `define AXI_B_LAYER_M3_S9 `i_axi_AXI_B_LAYER_M3_S9
`endif 

`ifdef i_axi_AXI_B_LAYER_M3_S10
  `define AXI_B_LAYER_M3_S10 `i_axi_AXI_B_LAYER_M3_S10
`endif 

`ifdef i_axi_AXI_B_LAYER_M3_S11
  `define AXI_B_LAYER_M3_S11 `i_axi_AXI_B_LAYER_M3_S11
`endif 

`ifdef i_axi_AXI_B_LAYER_M3_S12
  `define AXI_B_LAYER_M3_S12 `i_axi_AXI_B_LAYER_M3_S12
`endif 

`ifdef i_axi_AXI_B_LAYER_M3_S13
  `define AXI_B_LAYER_M3_S13 `i_axi_AXI_B_LAYER_M3_S13
`endif 

`ifdef i_axi_AXI_B_LAYER_M3_S14
  `define AXI_B_LAYER_M3_S14 `i_axi_AXI_B_LAYER_M3_S14
`endif 

`ifdef i_axi_AXI_B_LAYER_M3_S15
  `define AXI_B_LAYER_M3_S15 `i_axi_AXI_B_LAYER_M3_S15
`endif 

`ifdef i_axi_AXI_B_LAYER_M3_S16
  `define AXI_B_LAYER_M3_S16 `i_axi_AXI_B_LAYER_M3_S16
`endif 

`ifdef i_axi_AXI_R_LAYER_M4_S0
  `define AXI_R_LAYER_M4_S0 `i_axi_AXI_R_LAYER_M4_S0
`endif 

`ifdef i_axi_AXI_R_LAYER_M4_S1
  `define AXI_R_LAYER_M4_S1 `i_axi_AXI_R_LAYER_M4_S1
`endif 

`ifdef i_axi_AXI_R_LAYER_M4_S2
  `define AXI_R_LAYER_M4_S2 `i_axi_AXI_R_LAYER_M4_S2
`endif 

`ifdef i_axi_AXI_R_LAYER_M4_S3
  `define AXI_R_LAYER_M4_S3 `i_axi_AXI_R_LAYER_M4_S3
`endif 

`ifdef i_axi_AXI_R_LAYER_M4_S4
  `define AXI_R_LAYER_M4_S4 `i_axi_AXI_R_LAYER_M4_S4
`endif 

`ifdef i_axi_AXI_R_LAYER_M4_S5
  `define AXI_R_LAYER_M4_S5 `i_axi_AXI_R_LAYER_M4_S5
`endif 

`ifdef i_axi_AXI_R_LAYER_M4_S6
  `define AXI_R_LAYER_M4_S6 `i_axi_AXI_R_LAYER_M4_S6
`endif 

`ifdef i_axi_AXI_R_LAYER_M4_S7
  `define AXI_R_LAYER_M4_S7 `i_axi_AXI_R_LAYER_M4_S7
`endif 

`ifdef i_axi_AXI_R_LAYER_M4_S8
  `define AXI_R_LAYER_M4_S8 `i_axi_AXI_R_LAYER_M4_S8
`endif 

`ifdef i_axi_AXI_R_LAYER_M4_S9
  `define AXI_R_LAYER_M4_S9 `i_axi_AXI_R_LAYER_M4_S9
`endif 

`ifdef i_axi_AXI_R_LAYER_M4_S10
  `define AXI_R_LAYER_M4_S10 `i_axi_AXI_R_LAYER_M4_S10
`endif 

`ifdef i_axi_AXI_R_LAYER_M4_S11
  `define AXI_R_LAYER_M4_S11 `i_axi_AXI_R_LAYER_M4_S11
`endif 

`ifdef i_axi_AXI_R_LAYER_M4_S12
  `define AXI_R_LAYER_M4_S12 `i_axi_AXI_R_LAYER_M4_S12
`endif 

`ifdef i_axi_AXI_R_LAYER_M4_S13
  `define AXI_R_LAYER_M4_S13 `i_axi_AXI_R_LAYER_M4_S13
`endif 

`ifdef i_axi_AXI_R_LAYER_M4_S14
  `define AXI_R_LAYER_M4_S14 `i_axi_AXI_R_LAYER_M4_S14
`endif 

`ifdef i_axi_AXI_R_LAYER_M4_S15
  `define AXI_R_LAYER_M4_S15 `i_axi_AXI_R_LAYER_M4_S15
`endif 

`ifdef i_axi_AXI_R_LAYER_M4_S16
  `define AXI_R_LAYER_M4_S16 `i_axi_AXI_R_LAYER_M4_S16
`endif 

`ifdef i_axi_AXI_B_LAYER_M4_S0
  `define AXI_B_LAYER_M4_S0 `i_axi_AXI_B_LAYER_M4_S0
`endif 

`ifdef i_axi_AXI_B_LAYER_M4_S1
  `define AXI_B_LAYER_M4_S1 `i_axi_AXI_B_LAYER_M4_S1
`endif 

`ifdef i_axi_AXI_B_LAYER_M4_S2
  `define AXI_B_LAYER_M4_S2 `i_axi_AXI_B_LAYER_M4_S2
`endif 

`ifdef i_axi_AXI_B_LAYER_M4_S3
  `define AXI_B_LAYER_M4_S3 `i_axi_AXI_B_LAYER_M4_S3
`endif 

`ifdef i_axi_AXI_B_LAYER_M4_S4
  `define AXI_B_LAYER_M4_S4 `i_axi_AXI_B_LAYER_M4_S4
`endif 

`ifdef i_axi_AXI_B_LAYER_M4_S5
  `define AXI_B_LAYER_M4_S5 `i_axi_AXI_B_LAYER_M4_S5
`endif 

`ifdef i_axi_AXI_B_LAYER_M4_S6
  `define AXI_B_LAYER_M4_S6 `i_axi_AXI_B_LAYER_M4_S6
`endif 

`ifdef i_axi_AXI_B_LAYER_M4_S7
  `define AXI_B_LAYER_M4_S7 `i_axi_AXI_B_LAYER_M4_S7
`endif 

`ifdef i_axi_AXI_B_LAYER_M4_S8
  `define AXI_B_LAYER_M4_S8 `i_axi_AXI_B_LAYER_M4_S8
`endif 

`ifdef i_axi_AXI_B_LAYER_M4_S9
  `define AXI_B_LAYER_M4_S9 `i_axi_AXI_B_LAYER_M4_S9
`endif 

`ifdef i_axi_AXI_B_LAYER_M4_S10
  `define AXI_B_LAYER_M4_S10 `i_axi_AXI_B_LAYER_M4_S10
`endif 

`ifdef i_axi_AXI_B_LAYER_M4_S11
  `define AXI_B_LAYER_M4_S11 `i_axi_AXI_B_LAYER_M4_S11
`endif 

`ifdef i_axi_AXI_B_LAYER_M4_S12
  `define AXI_B_LAYER_M4_S12 `i_axi_AXI_B_LAYER_M4_S12
`endif 

`ifdef i_axi_AXI_B_LAYER_M4_S13
  `define AXI_B_LAYER_M4_S13 `i_axi_AXI_B_LAYER_M4_S13
`endif 

`ifdef i_axi_AXI_B_LAYER_M4_S14
  `define AXI_B_LAYER_M4_S14 `i_axi_AXI_B_LAYER_M4_S14
`endif 

`ifdef i_axi_AXI_B_LAYER_M4_S15
  `define AXI_B_LAYER_M4_S15 `i_axi_AXI_B_LAYER_M4_S15
`endif 

`ifdef i_axi_AXI_B_LAYER_M4_S16
  `define AXI_B_LAYER_M4_S16 `i_axi_AXI_B_LAYER_M4_S16
`endif 

`ifdef i_axi_AXI_R_LAYER_M5_S0
  `define AXI_R_LAYER_M5_S0 `i_axi_AXI_R_LAYER_M5_S0
`endif 

`ifdef i_axi_AXI_R_LAYER_M5_S1
  `define AXI_R_LAYER_M5_S1 `i_axi_AXI_R_LAYER_M5_S1
`endif 

`ifdef i_axi_AXI_R_LAYER_M5_S2
  `define AXI_R_LAYER_M5_S2 `i_axi_AXI_R_LAYER_M5_S2
`endif 

`ifdef i_axi_AXI_R_LAYER_M5_S3
  `define AXI_R_LAYER_M5_S3 `i_axi_AXI_R_LAYER_M5_S3
`endif 

`ifdef i_axi_AXI_R_LAYER_M5_S4
  `define AXI_R_LAYER_M5_S4 `i_axi_AXI_R_LAYER_M5_S4
`endif 

`ifdef i_axi_AXI_R_LAYER_M5_S5
  `define AXI_R_LAYER_M5_S5 `i_axi_AXI_R_LAYER_M5_S5
`endif 

`ifdef i_axi_AXI_R_LAYER_M5_S6
  `define AXI_R_LAYER_M5_S6 `i_axi_AXI_R_LAYER_M5_S6
`endif 

`ifdef i_axi_AXI_R_LAYER_M5_S7
  `define AXI_R_LAYER_M5_S7 `i_axi_AXI_R_LAYER_M5_S7
`endif 

`ifdef i_axi_AXI_R_LAYER_M5_S8
  `define AXI_R_LAYER_M5_S8 `i_axi_AXI_R_LAYER_M5_S8
`endif 

`ifdef i_axi_AXI_R_LAYER_M5_S9
  `define AXI_R_LAYER_M5_S9 `i_axi_AXI_R_LAYER_M5_S9
`endif 

`ifdef i_axi_AXI_R_LAYER_M5_S10
  `define AXI_R_LAYER_M5_S10 `i_axi_AXI_R_LAYER_M5_S10
`endif 

`ifdef i_axi_AXI_R_LAYER_M5_S11
  `define AXI_R_LAYER_M5_S11 `i_axi_AXI_R_LAYER_M5_S11
`endif 

`ifdef i_axi_AXI_R_LAYER_M5_S12
  `define AXI_R_LAYER_M5_S12 `i_axi_AXI_R_LAYER_M5_S12
`endif 

`ifdef i_axi_AXI_R_LAYER_M5_S13
  `define AXI_R_LAYER_M5_S13 `i_axi_AXI_R_LAYER_M5_S13
`endif 

`ifdef i_axi_AXI_R_LAYER_M5_S14
  `define AXI_R_LAYER_M5_S14 `i_axi_AXI_R_LAYER_M5_S14
`endif 

`ifdef i_axi_AXI_R_LAYER_M5_S15
  `define AXI_R_LAYER_M5_S15 `i_axi_AXI_R_LAYER_M5_S15
`endif 

`ifdef i_axi_AXI_R_LAYER_M5_S16
  `define AXI_R_LAYER_M5_S16 `i_axi_AXI_R_LAYER_M5_S16
`endif 

`ifdef i_axi_AXI_B_LAYER_M5_S0
  `define AXI_B_LAYER_M5_S0 `i_axi_AXI_B_LAYER_M5_S0
`endif 

`ifdef i_axi_AXI_B_LAYER_M5_S1
  `define AXI_B_LAYER_M5_S1 `i_axi_AXI_B_LAYER_M5_S1
`endif 

`ifdef i_axi_AXI_B_LAYER_M5_S2
  `define AXI_B_LAYER_M5_S2 `i_axi_AXI_B_LAYER_M5_S2
`endif 

`ifdef i_axi_AXI_B_LAYER_M5_S3
  `define AXI_B_LAYER_M5_S3 `i_axi_AXI_B_LAYER_M5_S3
`endif 

`ifdef i_axi_AXI_B_LAYER_M5_S4
  `define AXI_B_LAYER_M5_S4 `i_axi_AXI_B_LAYER_M5_S4
`endif 

`ifdef i_axi_AXI_B_LAYER_M5_S5
  `define AXI_B_LAYER_M5_S5 `i_axi_AXI_B_LAYER_M5_S5
`endif 

`ifdef i_axi_AXI_B_LAYER_M5_S6
  `define AXI_B_LAYER_M5_S6 `i_axi_AXI_B_LAYER_M5_S6
`endif 

`ifdef i_axi_AXI_B_LAYER_M5_S7
  `define AXI_B_LAYER_M5_S7 `i_axi_AXI_B_LAYER_M5_S7
`endif 

`ifdef i_axi_AXI_B_LAYER_M5_S8
  `define AXI_B_LAYER_M5_S8 `i_axi_AXI_B_LAYER_M5_S8
`endif 

`ifdef i_axi_AXI_B_LAYER_M5_S9
  `define AXI_B_LAYER_M5_S9 `i_axi_AXI_B_LAYER_M5_S9
`endif 

`ifdef i_axi_AXI_B_LAYER_M5_S10
  `define AXI_B_LAYER_M5_S10 `i_axi_AXI_B_LAYER_M5_S10
`endif 

`ifdef i_axi_AXI_B_LAYER_M5_S11
  `define AXI_B_LAYER_M5_S11 `i_axi_AXI_B_LAYER_M5_S11
`endif 

`ifdef i_axi_AXI_B_LAYER_M5_S12
  `define AXI_B_LAYER_M5_S12 `i_axi_AXI_B_LAYER_M5_S12
`endif 

`ifdef i_axi_AXI_B_LAYER_M5_S13
  `define AXI_B_LAYER_M5_S13 `i_axi_AXI_B_LAYER_M5_S13
`endif 

`ifdef i_axi_AXI_B_LAYER_M5_S14
  `define AXI_B_LAYER_M5_S14 `i_axi_AXI_B_LAYER_M5_S14
`endif 

`ifdef i_axi_AXI_B_LAYER_M5_S15
  `define AXI_B_LAYER_M5_S15 `i_axi_AXI_B_LAYER_M5_S15
`endif 

`ifdef i_axi_AXI_B_LAYER_M5_S16
  `define AXI_B_LAYER_M5_S16 `i_axi_AXI_B_LAYER_M5_S16
`endif 

`ifdef i_axi_AXI_R_LAYER_M6_S0
  `define AXI_R_LAYER_M6_S0 `i_axi_AXI_R_LAYER_M6_S0
`endif 

`ifdef i_axi_AXI_R_LAYER_M6_S1
  `define AXI_R_LAYER_M6_S1 `i_axi_AXI_R_LAYER_M6_S1
`endif 

`ifdef i_axi_AXI_R_LAYER_M6_S2
  `define AXI_R_LAYER_M6_S2 `i_axi_AXI_R_LAYER_M6_S2
`endif 

`ifdef i_axi_AXI_R_LAYER_M6_S3
  `define AXI_R_LAYER_M6_S3 `i_axi_AXI_R_LAYER_M6_S3
`endif 

`ifdef i_axi_AXI_R_LAYER_M6_S4
  `define AXI_R_LAYER_M6_S4 `i_axi_AXI_R_LAYER_M6_S4
`endif 

`ifdef i_axi_AXI_R_LAYER_M6_S5
  `define AXI_R_LAYER_M6_S5 `i_axi_AXI_R_LAYER_M6_S5
`endif 

`ifdef i_axi_AXI_R_LAYER_M6_S6
  `define AXI_R_LAYER_M6_S6 `i_axi_AXI_R_LAYER_M6_S6
`endif 

`ifdef i_axi_AXI_R_LAYER_M6_S7
  `define AXI_R_LAYER_M6_S7 `i_axi_AXI_R_LAYER_M6_S7
`endif 

`ifdef i_axi_AXI_R_LAYER_M6_S8
  `define AXI_R_LAYER_M6_S8 `i_axi_AXI_R_LAYER_M6_S8
`endif 

`ifdef i_axi_AXI_R_LAYER_M6_S9
  `define AXI_R_LAYER_M6_S9 `i_axi_AXI_R_LAYER_M6_S9
`endif 

`ifdef i_axi_AXI_R_LAYER_M6_S10
  `define AXI_R_LAYER_M6_S10 `i_axi_AXI_R_LAYER_M6_S10
`endif 

`ifdef i_axi_AXI_R_LAYER_M6_S11
  `define AXI_R_LAYER_M6_S11 `i_axi_AXI_R_LAYER_M6_S11
`endif 

`ifdef i_axi_AXI_R_LAYER_M6_S12
  `define AXI_R_LAYER_M6_S12 `i_axi_AXI_R_LAYER_M6_S12
`endif 

`ifdef i_axi_AXI_R_LAYER_M6_S13
  `define AXI_R_LAYER_M6_S13 `i_axi_AXI_R_LAYER_M6_S13
`endif 

`ifdef i_axi_AXI_R_LAYER_M6_S14
  `define AXI_R_LAYER_M6_S14 `i_axi_AXI_R_LAYER_M6_S14
`endif 

`ifdef i_axi_AXI_R_LAYER_M6_S15
  `define AXI_R_LAYER_M6_S15 `i_axi_AXI_R_LAYER_M6_S15
`endif 

`ifdef i_axi_AXI_R_LAYER_M6_S16
  `define AXI_R_LAYER_M6_S16 `i_axi_AXI_R_LAYER_M6_S16
`endif 

`ifdef i_axi_AXI_B_LAYER_M6_S0
  `define AXI_B_LAYER_M6_S0 `i_axi_AXI_B_LAYER_M6_S0
`endif 

`ifdef i_axi_AXI_B_LAYER_M6_S1
  `define AXI_B_LAYER_M6_S1 `i_axi_AXI_B_LAYER_M6_S1
`endif 

`ifdef i_axi_AXI_B_LAYER_M6_S2
  `define AXI_B_LAYER_M6_S2 `i_axi_AXI_B_LAYER_M6_S2
`endif 

`ifdef i_axi_AXI_B_LAYER_M6_S3
  `define AXI_B_LAYER_M6_S3 `i_axi_AXI_B_LAYER_M6_S3
`endif 

`ifdef i_axi_AXI_B_LAYER_M6_S4
  `define AXI_B_LAYER_M6_S4 `i_axi_AXI_B_LAYER_M6_S4
`endif 

`ifdef i_axi_AXI_B_LAYER_M6_S5
  `define AXI_B_LAYER_M6_S5 `i_axi_AXI_B_LAYER_M6_S5
`endif 

`ifdef i_axi_AXI_B_LAYER_M6_S6
  `define AXI_B_LAYER_M6_S6 `i_axi_AXI_B_LAYER_M6_S6
`endif 

`ifdef i_axi_AXI_B_LAYER_M6_S7
  `define AXI_B_LAYER_M6_S7 `i_axi_AXI_B_LAYER_M6_S7
`endif 

`ifdef i_axi_AXI_B_LAYER_M6_S8
  `define AXI_B_LAYER_M6_S8 `i_axi_AXI_B_LAYER_M6_S8
`endif 

`ifdef i_axi_AXI_B_LAYER_M6_S9
  `define AXI_B_LAYER_M6_S9 `i_axi_AXI_B_LAYER_M6_S9
`endif 

`ifdef i_axi_AXI_B_LAYER_M6_S10
  `define AXI_B_LAYER_M6_S10 `i_axi_AXI_B_LAYER_M6_S10
`endif 

`ifdef i_axi_AXI_B_LAYER_M6_S11
  `define AXI_B_LAYER_M6_S11 `i_axi_AXI_B_LAYER_M6_S11
`endif 

`ifdef i_axi_AXI_B_LAYER_M6_S12
  `define AXI_B_LAYER_M6_S12 `i_axi_AXI_B_LAYER_M6_S12
`endif 

`ifdef i_axi_AXI_B_LAYER_M6_S13
  `define AXI_B_LAYER_M6_S13 `i_axi_AXI_B_LAYER_M6_S13
`endif 

`ifdef i_axi_AXI_B_LAYER_M6_S14
  `define AXI_B_LAYER_M6_S14 `i_axi_AXI_B_LAYER_M6_S14
`endif 

`ifdef i_axi_AXI_B_LAYER_M6_S15
  `define AXI_B_LAYER_M6_S15 `i_axi_AXI_B_LAYER_M6_S15
`endif 

`ifdef i_axi_AXI_B_LAYER_M6_S16
  `define AXI_B_LAYER_M6_S16 `i_axi_AXI_B_LAYER_M6_S16
`endif 

`ifdef i_axi_AXI_R_LAYER_M7_S0
  `define AXI_R_LAYER_M7_S0 `i_axi_AXI_R_LAYER_M7_S0
`endif 

`ifdef i_axi_AXI_R_LAYER_M7_S1
  `define AXI_R_LAYER_M7_S1 `i_axi_AXI_R_LAYER_M7_S1
`endif 

`ifdef i_axi_AXI_R_LAYER_M7_S2
  `define AXI_R_LAYER_M7_S2 `i_axi_AXI_R_LAYER_M7_S2
`endif 

`ifdef i_axi_AXI_R_LAYER_M7_S3
  `define AXI_R_LAYER_M7_S3 `i_axi_AXI_R_LAYER_M7_S3
`endif 

`ifdef i_axi_AXI_R_LAYER_M7_S4
  `define AXI_R_LAYER_M7_S4 `i_axi_AXI_R_LAYER_M7_S4
`endif 

`ifdef i_axi_AXI_R_LAYER_M7_S5
  `define AXI_R_LAYER_M7_S5 `i_axi_AXI_R_LAYER_M7_S5
`endif 

`ifdef i_axi_AXI_R_LAYER_M7_S6
  `define AXI_R_LAYER_M7_S6 `i_axi_AXI_R_LAYER_M7_S6
`endif 

`ifdef i_axi_AXI_R_LAYER_M7_S7
  `define AXI_R_LAYER_M7_S7 `i_axi_AXI_R_LAYER_M7_S7
`endif 

`ifdef i_axi_AXI_R_LAYER_M7_S8
  `define AXI_R_LAYER_M7_S8 `i_axi_AXI_R_LAYER_M7_S8
`endif 

`ifdef i_axi_AXI_R_LAYER_M7_S9
  `define AXI_R_LAYER_M7_S9 `i_axi_AXI_R_LAYER_M7_S9
`endif 

`ifdef i_axi_AXI_R_LAYER_M7_S10
  `define AXI_R_LAYER_M7_S10 `i_axi_AXI_R_LAYER_M7_S10
`endif 

`ifdef i_axi_AXI_R_LAYER_M7_S11
  `define AXI_R_LAYER_M7_S11 `i_axi_AXI_R_LAYER_M7_S11
`endif 

`ifdef i_axi_AXI_R_LAYER_M7_S12
  `define AXI_R_LAYER_M7_S12 `i_axi_AXI_R_LAYER_M7_S12
`endif 

`ifdef i_axi_AXI_R_LAYER_M7_S13
  `define AXI_R_LAYER_M7_S13 `i_axi_AXI_R_LAYER_M7_S13
`endif 

`ifdef i_axi_AXI_R_LAYER_M7_S14
  `define AXI_R_LAYER_M7_S14 `i_axi_AXI_R_LAYER_M7_S14
`endif 

`ifdef i_axi_AXI_R_LAYER_M7_S15
  `define AXI_R_LAYER_M7_S15 `i_axi_AXI_R_LAYER_M7_S15
`endif 

`ifdef i_axi_AXI_R_LAYER_M7_S16
  `define AXI_R_LAYER_M7_S16 `i_axi_AXI_R_LAYER_M7_S16
`endif 

`ifdef i_axi_AXI_B_LAYER_M7_S0
  `define AXI_B_LAYER_M7_S0 `i_axi_AXI_B_LAYER_M7_S0
`endif 

`ifdef i_axi_AXI_B_LAYER_M7_S1
  `define AXI_B_LAYER_M7_S1 `i_axi_AXI_B_LAYER_M7_S1
`endif 

`ifdef i_axi_AXI_B_LAYER_M7_S2
  `define AXI_B_LAYER_M7_S2 `i_axi_AXI_B_LAYER_M7_S2
`endif 

`ifdef i_axi_AXI_B_LAYER_M7_S3
  `define AXI_B_LAYER_M7_S3 `i_axi_AXI_B_LAYER_M7_S3
`endif 

`ifdef i_axi_AXI_B_LAYER_M7_S4
  `define AXI_B_LAYER_M7_S4 `i_axi_AXI_B_LAYER_M7_S4
`endif 

`ifdef i_axi_AXI_B_LAYER_M7_S5
  `define AXI_B_LAYER_M7_S5 `i_axi_AXI_B_LAYER_M7_S5
`endif 

`ifdef i_axi_AXI_B_LAYER_M7_S6
  `define AXI_B_LAYER_M7_S6 `i_axi_AXI_B_LAYER_M7_S6
`endif 

`ifdef i_axi_AXI_B_LAYER_M7_S7
  `define AXI_B_LAYER_M7_S7 `i_axi_AXI_B_LAYER_M7_S7
`endif 

`ifdef i_axi_AXI_B_LAYER_M7_S8
  `define AXI_B_LAYER_M7_S8 `i_axi_AXI_B_LAYER_M7_S8
`endif 

`ifdef i_axi_AXI_B_LAYER_M7_S9
  `define AXI_B_LAYER_M7_S9 `i_axi_AXI_B_LAYER_M7_S9
`endif 

`ifdef i_axi_AXI_B_LAYER_M7_S10
  `define AXI_B_LAYER_M7_S10 `i_axi_AXI_B_LAYER_M7_S10
`endif 

`ifdef i_axi_AXI_B_LAYER_M7_S11
  `define AXI_B_LAYER_M7_S11 `i_axi_AXI_B_LAYER_M7_S11
`endif 

`ifdef i_axi_AXI_B_LAYER_M7_S12
  `define AXI_B_LAYER_M7_S12 `i_axi_AXI_B_LAYER_M7_S12
`endif 

`ifdef i_axi_AXI_B_LAYER_M7_S13
  `define AXI_B_LAYER_M7_S13 `i_axi_AXI_B_LAYER_M7_S13
`endif 

`ifdef i_axi_AXI_B_LAYER_M7_S14
  `define AXI_B_LAYER_M7_S14 `i_axi_AXI_B_LAYER_M7_S14
`endif 

`ifdef i_axi_AXI_B_LAYER_M7_S15
  `define AXI_B_LAYER_M7_S15 `i_axi_AXI_B_LAYER_M7_S15
`endif 

`ifdef i_axi_AXI_B_LAYER_M7_S16
  `define AXI_B_LAYER_M7_S16 `i_axi_AXI_B_LAYER_M7_S16
`endif 

`ifdef i_axi_AXI_R_LAYER_M8_S0
  `define AXI_R_LAYER_M8_S0 `i_axi_AXI_R_LAYER_M8_S0
`endif 

`ifdef i_axi_AXI_R_LAYER_M8_S1
  `define AXI_R_LAYER_M8_S1 `i_axi_AXI_R_LAYER_M8_S1
`endif 

`ifdef i_axi_AXI_R_LAYER_M8_S2
  `define AXI_R_LAYER_M8_S2 `i_axi_AXI_R_LAYER_M8_S2
`endif 

`ifdef i_axi_AXI_R_LAYER_M8_S3
  `define AXI_R_LAYER_M8_S3 `i_axi_AXI_R_LAYER_M8_S3
`endif 

`ifdef i_axi_AXI_R_LAYER_M8_S4
  `define AXI_R_LAYER_M8_S4 `i_axi_AXI_R_LAYER_M8_S4
`endif 

`ifdef i_axi_AXI_R_LAYER_M8_S5
  `define AXI_R_LAYER_M8_S5 `i_axi_AXI_R_LAYER_M8_S5
`endif 

`ifdef i_axi_AXI_R_LAYER_M8_S6
  `define AXI_R_LAYER_M8_S6 `i_axi_AXI_R_LAYER_M8_S6
`endif 

`ifdef i_axi_AXI_R_LAYER_M8_S7
  `define AXI_R_LAYER_M8_S7 `i_axi_AXI_R_LAYER_M8_S7
`endif 

`ifdef i_axi_AXI_R_LAYER_M8_S8
  `define AXI_R_LAYER_M8_S8 `i_axi_AXI_R_LAYER_M8_S8
`endif 

`ifdef i_axi_AXI_R_LAYER_M8_S9
  `define AXI_R_LAYER_M8_S9 `i_axi_AXI_R_LAYER_M8_S9
`endif 

`ifdef i_axi_AXI_R_LAYER_M8_S10
  `define AXI_R_LAYER_M8_S10 `i_axi_AXI_R_LAYER_M8_S10
`endif 

`ifdef i_axi_AXI_R_LAYER_M8_S11
  `define AXI_R_LAYER_M8_S11 `i_axi_AXI_R_LAYER_M8_S11
`endif 

`ifdef i_axi_AXI_R_LAYER_M8_S12
  `define AXI_R_LAYER_M8_S12 `i_axi_AXI_R_LAYER_M8_S12
`endif 

`ifdef i_axi_AXI_R_LAYER_M8_S13
  `define AXI_R_LAYER_M8_S13 `i_axi_AXI_R_LAYER_M8_S13
`endif 

`ifdef i_axi_AXI_R_LAYER_M8_S14
  `define AXI_R_LAYER_M8_S14 `i_axi_AXI_R_LAYER_M8_S14
`endif 

`ifdef i_axi_AXI_R_LAYER_M8_S15
  `define AXI_R_LAYER_M8_S15 `i_axi_AXI_R_LAYER_M8_S15
`endif 

`ifdef i_axi_AXI_R_LAYER_M8_S16
  `define AXI_R_LAYER_M8_S16 `i_axi_AXI_R_LAYER_M8_S16
`endif 

`ifdef i_axi_AXI_B_LAYER_M8_S0
  `define AXI_B_LAYER_M8_S0 `i_axi_AXI_B_LAYER_M8_S0
`endif 

`ifdef i_axi_AXI_B_LAYER_M8_S1
  `define AXI_B_LAYER_M8_S1 `i_axi_AXI_B_LAYER_M8_S1
`endif 

`ifdef i_axi_AXI_B_LAYER_M8_S2
  `define AXI_B_LAYER_M8_S2 `i_axi_AXI_B_LAYER_M8_S2
`endif 

`ifdef i_axi_AXI_B_LAYER_M8_S3
  `define AXI_B_LAYER_M8_S3 `i_axi_AXI_B_LAYER_M8_S3
`endif 

`ifdef i_axi_AXI_B_LAYER_M8_S4
  `define AXI_B_LAYER_M8_S4 `i_axi_AXI_B_LAYER_M8_S4
`endif 

`ifdef i_axi_AXI_B_LAYER_M8_S5
  `define AXI_B_LAYER_M8_S5 `i_axi_AXI_B_LAYER_M8_S5
`endif 

`ifdef i_axi_AXI_B_LAYER_M8_S6
  `define AXI_B_LAYER_M8_S6 `i_axi_AXI_B_LAYER_M8_S6
`endif 

`ifdef i_axi_AXI_B_LAYER_M8_S7
  `define AXI_B_LAYER_M8_S7 `i_axi_AXI_B_LAYER_M8_S7
`endif 

`ifdef i_axi_AXI_B_LAYER_M8_S8
  `define AXI_B_LAYER_M8_S8 `i_axi_AXI_B_LAYER_M8_S8
`endif 

`ifdef i_axi_AXI_B_LAYER_M8_S9
  `define AXI_B_LAYER_M8_S9 `i_axi_AXI_B_LAYER_M8_S9
`endif 

`ifdef i_axi_AXI_B_LAYER_M8_S10
  `define AXI_B_LAYER_M8_S10 `i_axi_AXI_B_LAYER_M8_S10
`endif 

`ifdef i_axi_AXI_B_LAYER_M8_S11
  `define AXI_B_LAYER_M8_S11 `i_axi_AXI_B_LAYER_M8_S11
`endif 

`ifdef i_axi_AXI_B_LAYER_M8_S12
  `define AXI_B_LAYER_M8_S12 `i_axi_AXI_B_LAYER_M8_S12
`endif 

`ifdef i_axi_AXI_B_LAYER_M8_S13
  `define AXI_B_LAYER_M8_S13 `i_axi_AXI_B_LAYER_M8_S13
`endif 

`ifdef i_axi_AXI_B_LAYER_M8_S14
  `define AXI_B_LAYER_M8_S14 `i_axi_AXI_B_LAYER_M8_S14
`endif 

`ifdef i_axi_AXI_B_LAYER_M8_S15
  `define AXI_B_LAYER_M8_S15 `i_axi_AXI_B_LAYER_M8_S15
`endif 

`ifdef i_axi_AXI_B_LAYER_M8_S16
  `define AXI_B_LAYER_M8_S16 `i_axi_AXI_B_LAYER_M8_S16
`endif 

`ifdef i_axi_AXI_R_LAYER_M9_S0
  `define AXI_R_LAYER_M9_S0 `i_axi_AXI_R_LAYER_M9_S0
`endif 

`ifdef i_axi_AXI_R_LAYER_M9_S1
  `define AXI_R_LAYER_M9_S1 `i_axi_AXI_R_LAYER_M9_S1
`endif 

`ifdef i_axi_AXI_R_LAYER_M9_S2
  `define AXI_R_LAYER_M9_S2 `i_axi_AXI_R_LAYER_M9_S2
`endif 

`ifdef i_axi_AXI_R_LAYER_M9_S3
  `define AXI_R_LAYER_M9_S3 `i_axi_AXI_R_LAYER_M9_S3
`endif 

`ifdef i_axi_AXI_R_LAYER_M9_S4
  `define AXI_R_LAYER_M9_S4 `i_axi_AXI_R_LAYER_M9_S4
`endif 

`ifdef i_axi_AXI_R_LAYER_M9_S5
  `define AXI_R_LAYER_M9_S5 `i_axi_AXI_R_LAYER_M9_S5
`endif 

`ifdef i_axi_AXI_R_LAYER_M9_S6
  `define AXI_R_LAYER_M9_S6 `i_axi_AXI_R_LAYER_M9_S6
`endif 

`ifdef i_axi_AXI_R_LAYER_M9_S7
  `define AXI_R_LAYER_M9_S7 `i_axi_AXI_R_LAYER_M9_S7
`endif 

`ifdef i_axi_AXI_R_LAYER_M9_S8
  `define AXI_R_LAYER_M9_S8 `i_axi_AXI_R_LAYER_M9_S8
`endif 

`ifdef i_axi_AXI_R_LAYER_M9_S9
  `define AXI_R_LAYER_M9_S9 `i_axi_AXI_R_LAYER_M9_S9
`endif 

`ifdef i_axi_AXI_R_LAYER_M9_S10
  `define AXI_R_LAYER_M9_S10 `i_axi_AXI_R_LAYER_M9_S10
`endif 

`ifdef i_axi_AXI_R_LAYER_M9_S11
  `define AXI_R_LAYER_M9_S11 `i_axi_AXI_R_LAYER_M9_S11
`endif 

`ifdef i_axi_AXI_R_LAYER_M9_S12
  `define AXI_R_LAYER_M9_S12 `i_axi_AXI_R_LAYER_M9_S12
`endif 

`ifdef i_axi_AXI_R_LAYER_M9_S13
  `define AXI_R_LAYER_M9_S13 `i_axi_AXI_R_LAYER_M9_S13
`endif 

`ifdef i_axi_AXI_R_LAYER_M9_S14
  `define AXI_R_LAYER_M9_S14 `i_axi_AXI_R_LAYER_M9_S14
`endif 

`ifdef i_axi_AXI_R_LAYER_M9_S15
  `define AXI_R_LAYER_M9_S15 `i_axi_AXI_R_LAYER_M9_S15
`endif 

`ifdef i_axi_AXI_R_LAYER_M9_S16
  `define AXI_R_LAYER_M9_S16 `i_axi_AXI_R_LAYER_M9_S16
`endif 

`ifdef i_axi_AXI_B_LAYER_M9_S0
  `define AXI_B_LAYER_M9_S0 `i_axi_AXI_B_LAYER_M9_S0
`endif 

`ifdef i_axi_AXI_B_LAYER_M9_S1
  `define AXI_B_LAYER_M9_S1 `i_axi_AXI_B_LAYER_M9_S1
`endif 

`ifdef i_axi_AXI_B_LAYER_M9_S2
  `define AXI_B_LAYER_M9_S2 `i_axi_AXI_B_LAYER_M9_S2
`endif 

`ifdef i_axi_AXI_B_LAYER_M9_S3
  `define AXI_B_LAYER_M9_S3 `i_axi_AXI_B_LAYER_M9_S3
`endif 

`ifdef i_axi_AXI_B_LAYER_M9_S4
  `define AXI_B_LAYER_M9_S4 `i_axi_AXI_B_LAYER_M9_S4
`endif 

`ifdef i_axi_AXI_B_LAYER_M9_S5
  `define AXI_B_LAYER_M9_S5 `i_axi_AXI_B_LAYER_M9_S5
`endif 

`ifdef i_axi_AXI_B_LAYER_M9_S6
  `define AXI_B_LAYER_M9_S6 `i_axi_AXI_B_LAYER_M9_S6
`endif 

`ifdef i_axi_AXI_B_LAYER_M9_S7
  `define AXI_B_LAYER_M9_S7 `i_axi_AXI_B_LAYER_M9_S7
`endif 

`ifdef i_axi_AXI_B_LAYER_M9_S8
  `define AXI_B_LAYER_M9_S8 `i_axi_AXI_B_LAYER_M9_S8
`endif 

`ifdef i_axi_AXI_B_LAYER_M9_S9
  `define AXI_B_LAYER_M9_S9 `i_axi_AXI_B_LAYER_M9_S9
`endif 

`ifdef i_axi_AXI_B_LAYER_M9_S10
  `define AXI_B_LAYER_M9_S10 `i_axi_AXI_B_LAYER_M9_S10
`endif 

`ifdef i_axi_AXI_B_LAYER_M9_S11
  `define AXI_B_LAYER_M9_S11 `i_axi_AXI_B_LAYER_M9_S11
`endif 

`ifdef i_axi_AXI_B_LAYER_M9_S12
  `define AXI_B_LAYER_M9_S12 `i_axi_AXI_B_LAYER_M9_S12
`endif 

`ifdef i_axi_AXI_B_LAYER_M9_S13
  `define AXI_B_LAYER_M9_S13 `i_axi_AXI_B_LAYER_M9_S13
`endif 

`ifdef i_axi_AXI_B_LAYER_M9_S14
  `define AXI_B_LAYER_M9_S14 `i_axi_AXI_B_LAYER_M9_S14
`endif 

`ifdef i_axi_AXI_B_LAYER_M9_S15
  `define AXI_B_LAYER_M9_S15 `i_axi_AXI_B_LAYER_M9_S15
`endif 

`ifdef i_axi_AXI_B_LAYER_M9_S16
  `define AXI_B_LAYER_M9_S16 `i_axi_AXI_B_LAYER_M9_S16
`endif 

`ifdef i_axi_AXI_R_LAYER_M10_S0
  `define AXI_R_LAYER_M10_S0 `i_axi_AXI_R_LAYER_M10_S0
`endif 

`ifdef i_axi_AXI_R_LAYER_M10_S1
  `define AXI_R_LAYER_M10_S1 `i_axi_AXI_R_LAYER_M10_S1
`endif 

`ifdef i_axi_AXI_R_LAYER_M10_S2
  `define AXI_R_LAYER_M10_S2 `i_axi_AXI_R_LAYER_M10_S2
`endif 

`ifdef i_axi_AXI_R_LAYER_M10_S3
  `define AXI_R_LAYER_M10_S3 `i_axi_AXI_R_LAYER_M10_S3
`endif 

`ifdef i_axi_AXI_R_LAYER_M10_S4
  `define AXI_R_LAYER_M10_S4 `i_axi_AXI_R_LAYER_M10_S4
`endif 

`ifdef i_axi_AXI_R_LAYER_M10_S5
  `define AXI_R_LAYER_M10_S5 `i_axi_AXI_R_LAYER_M10_S5
`endif 

`ifdef i_axi_AXI_R_LAYER_M10_S6
  `define AXI_R_LAYER_M10_S6 `i_axi_AXI_R_LAYER_M10_S6
`endif 

`ifdef i_axi_AXI_R_LAYER_M10_S7
  `define AXI_R_LAYER_M10_S7 `i_axi_AXI_R_LAYER_M10_S7
`endif 

`ifdef i_axi_AXI_R_LAYER_M10_S8
  `define AXI_R_LAYER_M10_S8 `i_axi_AXI_R_LAYER_M10_S8
`endif 

`ifdef i_axi_AXI_R_LAYER_M10_S9
  `define AXI_R_LAYER_M10_S9 `i_axi_AXI_R_LAYER_M10_S9
`endif 

`ifdef i_axi_AXI_R_LAYER_M10_S10
  `define AXI_R_LAYER_M10_S10 `i_axi_AXI_R_LAYER_M10_S10
`endif 

`ifdef i_axi_AXI_R_LAYER_M10_S11
  `define AXI_R_LAYER_M10_S11 `i_axi_AXI_R_LAYER_M10_S11
`endif 

`ifdef i_axi_AXI_R_LAYER_M10_S12
  `define AXI_R_LAYER_M10_S12 `i_axi_AXI_R_LAYER_M10_S12
`endif 

`ifdef i_axi_AXI_R_LAYER_M10_S13
  `define AXI_R_LAYER_M10_S13 `i_axi_AXI_R_LAYER_M10_S13
`endif 

`ifdef i_axi_AXI_R_LAYER_M10_S14
  `define AXI_R_LAYER_M10_S14 `i_axi_AXI_R_LAYER_M10_S14
`endif 

`ifdef i_axi_AXI_R_LAYER_M10_S15
  `define AXI_R_LAYER_M10_S15 `i_axi_AXI_R_LAYER_M10_S15
`endif 

`ifdef i_axi_AXI_R_LAYER_M10_S16
  `define AXI_R_LAYER_M10_S16 `i_axi_AXI_R_LAYER_M10_S16
`endif 

`ifdef i_axi_AXI_B_LAYER_M10_S0
  `define AXI_B_LAYER_M10_S0 `i_axi_AXI_B_LAYER_M10_S0
`endif 

`ifdef i_axi_AXI_B_LAYER_M10_S1
  `define AXI_B_LAYER_M10_S1 `i_axi_AXI_B_LAYER_M10_S1
`endif 

`ifdef i_axi_AXI_B_LAYER_M10_S2
  `define AXI_B_LAYER_M10_S2 `i_axi_AXI_B_LAYER_M10_S2
`endif 

`ifdef i_axi_AXI_B_LAYER_M10_S3
  `define AXI_B_LAYER_M10_S3 `i_axi_AXI_B_LAYER_M10_S3
`endif 

`ifdef i_axi_AXI_B_LAYER_M10_S4
  `define AXI_B_LAYER_M10_S4 `i_axi_AXI_B_LAYER_M10_S4
`endif 

`ifdef i_axi_AXI_B_LAYER_M10_S5
  `define AXI_B_LAYER_M10_S5 `i_axi_AXI_B_LAYER_M10_S5
`endif 

`ifdef i_axi_AXI_B_LAYER_M10_S6
  `define AXI_B_LAYER_M10_S6 `i_axi_AXI_B_LAYER_M10_S6
`endif 

`ifdef i_axi_AXI_B_LAYER_M10_S7
  `define AXI_B_LAYER_M10_S7 `i_axi_AXI_B_LAYER_M10_S7
`endif 

`ifdef i_axi_AXI_B_LAYER_M10_S8
  `define AXI_B_LAYER_M10_S8 `i_axi_AXI_B_LAYER_M10_S8
`endif 

`ifdef i_axi_AXI_B_LAYER_M10_S9
  `define AXI_B_LAYER_M10_S9 `i_axi_AXI_B_LAYER_M10_S9
`endif 

`ifdef i_axi_AXI_B_LAYER_M10_S10
  `define AXI_B_LAYER_M10_S10 `i_axi_AXI_B_LAYER_M10_S10
`endif 

`ifdef i_axi_AXI_B_LAYER_M10_S11
  `define AXI_B_LAYER_M10_S11 `i_axi_AXI_B_LAYER_M10_S11
`endif 

`ifdef i_axi_AXI_B_LAYER_M10_S12
  `define AXI_B_LAYER_M10_S12 `i_axi_AXI_B_LAYER_M10_S12
`endif 

`ifdef i_axi_AXI_B_LAYER_M10_S13
  `define AXI_B_LAYER_M10_S13 `i_axi_AXI_B_LAYER_M10_S13
`endif 

`ifdef i_axi_AXI_B_LAYER_M10_S14
  `define AXI_B_LAYER_M10_S14 `i_axi_AXI_B_LAYER_M10_S14
`endif 

`ifdef i_axi_AXI_B_LAYER_M10_S15
  `define AXI_B_LAYER_M10_S15 `i_axi_AXI_B_LAYER_M10_S15
`endif 

`ifdef i_axi_AXI_B_LAYER_M10_S16
  `define AXI_B_LAYER_M10_S16 `i_axi_AXI_B_LAYER_M10_S16
`endif 

`ifdef i_axi_AXI_R_LAYER_M11_S0
  `define AXI_R_LAYER_M11_S0 `i_axi_AXI_R_LAYER_M11_S0
`endif 

`ifdef i_axi_AXI_R_LAYER_M11_S1
  `define AXI_R_LAYER_M11_S1 `i_axi_AXI_R_LAYER_M11_S1
`endif 

`ifdef i_axi_AXI_R_LAYER_M11_S2
  `define AXI_R_LAYER_M11_S2 `i_axi_AXI_R_LAYER_M11_S2
`endif 

`ifdef i_axi_AXI_R_LAYER_M11_S3
  `define AXI_R_LAYER_M11_S3 `i_axi_AXI_R_LAYER_M11_S3
`endif 

`ifdef i_axi_AXI_R_LAYER_M11_S4
  `define AXI_R_LAYER_M11_S4 `i_axi_AXI_R_LAYER_M11_S4
`endif 

`ifdef i_axi_AXI_R_LAYER_M11_S5
  `define AXI_R_LAYER_M11_S5 `i_axi_AXI_R_LAYER_M11_S5
`endif 

`ifdef i_axi_AXI_R_LAYER_M11_S6
  `define AXI_R_LAYER_M11_S6 `i_axi_AXI_R_LAYER_M11_S6
`endif 

`ifdef i_axi_AXI_R_LAYER_M11_S7
  `define AXI_R_LAYER_M11_S7 `i_axi_AXI_R_LAYER_M11_S7
`endif 

`ifdef i_axi_AXI_R_LAYER_M11_S8
  `define AXI_R_LAYER_M11_S8 `i_axi_AXI_R_LAYER_M11_S8
`endif 

`ifdef i_axi_AXI_R_LAYER_M11_S9
  `define AXI_R_LAYER_M11_S9 `i_axi_AXI_R_LAYER_M11_S9
`endif 

`ifdef i_axi_AXI_R_LAYER_M11_S10
  `define AXI_R_LAYER_M11_S10 `i_axi_AXI_R_LAYER_M11_S10
`endif 

`ifdef i_axi_AXI_R_LAYER_M11_S11
  `define AXI_R_LAYER_M11_S11 `i_axi_AXI_R_LAYER_M11_S11
`endif 

`ifdef i_axi_AXI_R_LAYER_M11_S12
  `define AXI_R_LAYER_M11_S12 `i_axi_AXI_R_LAYER_M11_S12
`endif 

`ifdef i_axi_AXI_R_LAYER_M11_S13
  `define AXI_R_LAYER_M11_S13 `i_axi_AXI_R_LAYER_M11_S13
`endif 

`ifdef i_axi_AXI_R_LAYER_M11_S14
  `define AXI_R_LAYER_M11_S14 `i_axi_AXI_R_LAYER_M11_S14
`endif 

`ifdef i_axi_AXI_R_LAYER_M11_S15
  `define AXI_R_LAYER_M11_S15 `i_axi_AXI_R_LAYER_M11_S15
`endif 

`ifdef i_axi_AXI_R_LAYER_M11_S16
  `define AXI_R_LAYER_M11_S16 `i_axi_AXI_R_LAYER_M11_S16
`endif 

`ifdef i_axi_AXI_B_LAYER_M11_S0
  `define AXI_B_LAYER_M11_S0 `i_axi_AXI_B_LAYER_M11_S0
`endif 

`ifdef i_axi_AXI_B_LAYER_M11_S1
  `define AXI_B_LAYER_M11_S1 `i_axi_AXI_B_LAYER_M11_S1
`endif 

`ifdef i_axi_AXI_B_LAYER_M11_S2
  `define AXI_B_LAYER_M11_S2 `i_axi_AXI_B_LAYER_M11_S2
`endif 

`ifdef i_axi_AXI_B_LAYER_M11_S3
  `define AXI_B_LAYER_M11_S3 `i_axi_AXI_B_LAYER_M11_S3
`endif 

`ifdef i_axi_AXI_B_LAYER_M11_S4
  `define AXI_B_LAYER_M11_S4 `i_axi_AXI_B_LAYER_M11_S4
`endif 

`ifdef i_axi_AXI_B_LAYER_M11_S5
  `define AXI_B_LAYER_M11_S5 `i_axi_AXI_B_LAYER_M11_S5
`endif 

`ifdef i_axi_AXI_B_LAYER_M11_S6
  `define AXI_B_LAYER_M11_S6 `i_axi_AXI_B_LAYER_M11_S6
`endif 

`ifdef i_axi_AXI_B_LAYER_M11_S7
  `define AXI_B_LAYER_M11_S7 `i_axi_AXI_B_LAYER_M11_S7
`endif 

`ifdef i_axi_AXI_B_LAYER_M11_S8
  `define AXI_B_LAYER_M11_S8 `i_axi_AXI_B_LAYER_M11_S8
`endif 

`ifdef i_axi_AXI_B_LAYER_M11_S9
  `define AXI_B_LAYER_M11_S9 `i_axi_AXI_B_LAYER_M11_S9
`endif 

`ifdef i_axi_AXI_B_LAYER_M11_S10
  `define AXI_B_LAYER_M11_S10 `i_axi_AXI_B_LAYER_M11_S10
`endif 

`ifdef i_axi_AXI_B_LAYER_M11_S11
  `define AXI_B_LAYER_M11_S11 `i_axi_AXI_B_LAYER_M11_S11
`endif 

`ifdef i_axi_AXI_B_LAYER_M11_S12
  `define AXI_B_LAYER_M11_S12 `i_axi_AXI_B_LAYER_M11_S12
`endif 

`ifdef i_axi_AXI_B_LAYER_M11_S13
  `define AXI_B_LAYER_M11_S13 `i_axi_AXI_B_LAYER_M11_S13
`endif 

`ifdef i_axi_AXI_B_LAYER_M11_S14
  `define AXI_B_LAYER_M11_S14 `i_axi_AXI_B_LAYER_M11_S14
`endif 

`ifdef i_axi_AXI_B_LAYER_M11_S15
  `define AXI_B_LAYER_M11_S15 `i_axi_AXI_B_LAYER_M11_S15
`endif 

`ifdef i_axi_AXI_B_LAYER_M11_S16
  `define AXI_B_LAYER_M11_S16 `i_axi_AXI_B_LAYER_M11_S16
`endif 

`ifdef i_axi_AXI_R_LAYER_M12_S0
  `define AXI_R_LAYER_M12_S0 `i_axi_AXI_R_LAYER_M12_S0
`endif 

`ifdef i_axi_AXI_R_LAYER_M12_S1
  `define AXI_R_LAYER_M12_S1 `i_axi_AXI_R_LAYER_M12_S1
`endif 

`ifdef i_axi_AXI_R_LAYER_M12_S2
  `define AXI_R_LAYER_M12_S2 `i_axi_AXI_R_LAYER_M12_S2
`endif 

`ifdef i_axi_AXI_R_LAYER_M12_S3
  `define AXI_R_LAYER_M12_S3 `i_axi_AXI_R_LAYER_M12_S3
`endif 

`ifdef i_axi_AXI_R_LAYER_M12_S4
  `define AXI_R_LAYER_M12_S4 `i_axi_AXI_R_LAYER_M12_S4
`endif 

`ifdef i_axi_AXI_R_LAYER_M12_S5
  `define AXI_R_LAYER_M12_S5 `i_axi_AXI_R_LAYER_M12_S5
`endif 

`ifdef i_axi_AXI_R_LAYER_M12_S6
  `define AXI_R_LAYER_M12_S6 `i_axi_AXI_R_LAYER_M12_S6
`endif 

`ifdef i_axi_AXI_R_LAYER_M12_S7
  `define AXI_R_LAYER_M12_S7 `i_axi_AXI_R_LAYER_M12_S7
`endif 

`ifdef i_axi_AXI_R_LAYER_M12_S8
  `define AXI_R_LAYER_M12_S8 `i_axi_AXI_R_LAYER_M12_S8
`endif 

`ifdef i_axi_AXI_R_LAYER_M12_S9
  `define AXI_R_LAYER_M12_S9 `i_axi_AXI_R_LAYER_M12_S9
`endif 

`ifdef i_axi_AXI_R_LAYER_M12_S10
  `define AXI_R_LAYER_M12_S10 `i_axi_AXI_R_LAYER_M12_S10
`endif 

`ifdef i_axi_AXI_R_LAYER_M12_S11
  `define AXI_R_LAYER_M12_S11 `i_axi_AXI_R_LAYER_M12_S11
`endif 

`ifdef i_axi_AXI_R_LAYER_M12_S12
  `define AXI_R_LAYER_M12_S12 `i_axi_AXI_R_LAYER_M12_S12
`endif 

`ifdef i_axi_AXI_R_LAYER_M12_S13
  `define AXI_R_LAYER_M12_S13 `i_axi_AXI_R_LAYER_M12_S13
`endif 

`ifdef i_axi_AXI_R_LAYER_M12_S14
  `define AXI_R_LAYER_M12_S14 `i_axi_AXI_R_LAYER_M12_S14
`endif 

`ifdef i_axi_AXI_R_LAYER_M12_S15
  `define AXI_R_LAYER_M12_S15 `i_axi_AXI_R_LAYER_M12_S15
`endif 

`ifdef i_axi_AXI_R_LAYER_M12_S16
  `define AXI_R_LAYER_M12_S16 `i_axi_AXI_R_LAYER_M12_S16
`endif 

`ifdef i_axi_AXI_B_LAYER_M12_S0
  `define AXI_B_LAYER_M12_S0 `i_axi_AXI_B_LAYER_M12_S0
`endif 

`ifdef i_axi_AXI_B_LAYER_M12_S1
  `define AXI_B_LAYER_M12_S1 `i_axi_AXI_B_LAYER_M12_S1
`endif 

`ifdef i_axi_AXI_B_LAYER_M12_S2
  `define AXI_B_LAYER_M12_S2 `i_axi_AXI_B_LAYER_M12_S2
`endif 

`ifdef i_axi_AXI_B_LAYER_M12_S3
  `define AXI_B_LAYER_M12_S3 `i_axi_AXI_B_LAYER_M12_S3
`endif 

`ifdef i_axi_AXI_B_LAYER_M12_S4
  `define AXI_B_LAYER_M12_S4 `i_axi_AXI_B_LAYER_M12_S4
`endif 

`ifdef i_axi_AXI_B_LAYER_M12_S5
  `define AXI_B_LAYER_M12_S5 `i_axi_AXI_B_LAYER_M12_S5
`endif 

`ifdef i_axi_AXI_B_LAYER_M12_S6
  `define AXI_B_LAYER_M12_S6 `i_axi_AXI_B_LAYER_M12_S6
`endif 

`ifdef i_axi_AXI_B_LAYER_M12_S7
  `define AXI_B_LAYER_M12_S7 `i_axi_AXI_B_LAYER_M12_S7
`endif 

`ifdef i_axi_AXI_B_LAYER_M12_S8
  `define AXI_B_LAYER_M12_S8 `i_axi_AXI_B_LAYER_M12_S8
`endif 

`ifdef i_axi_AXI_B_LAYER_M12_S9
  `define AXI_B_LAYER_M12_S9 `i_axi_AXI_B_LAYER_M12_S9
`endif 

`ifdef i_axi_AXI_B_LAYER_M12_S10
  `define AXI_B_LAYER_M12_S10 `i_axi_AXI_B_LAYER_M12_S10
`endif 

`ifdef i_axi_AXI_B_LAYER_M12_S11
  `define AXI_B_LAYER_M12_S11 `i_axi_AXI_B_LAYER_M12_S11
`endif 

`ifdef i_axi_AXI_B_LAYER_M12_S12
  `define AXI_B_LAYER_M12_S12 `i_axi_AXI_B_LAYER_M12_S12
`endif 

`ifdef i_axi_AXI_B_LAYER_M12_S13
  `define AXI_B_LAYER_M12_S13 `i_axi_AXI_B_LAYER_M12_S13
`endif 

`ifdef i_axi_AXI_B_LAYER_M12_S14
  `define AXI_B_LAYER_M12_S14 `i_axi_AXI_B_LAYER_M12_S14
`endif 

`ifdef i_axi_AXI_B_LAYER_M12_S15
  `define AXI_B_LAYER_M12_S15 `i_axi_AXI_B_LAYER_M12_S15
`endif 

`ifdef i_axi_AXI_B_LAYER_M12_S16
  `define AXI_B_LAYER_M12_S16 `i_axi_AXI_B_LAYER_M12_S16
`endif 

`ifdef i_axi_AXI_R_LAYER_M13_S0
  `define AXI_R_LAYER_M13_S0 `i_axi_AXI_R_LAYER_M13_S0
`endif 

`ifdef i_axi_AXI_R_LAYER_M13_S1
  `define AXI_R_LAYER_M13_S1 `i_axi_AXI_R_LAYER_M13_S1
`endif 

`ifdef i_axi_AXI_R_LAYER_M13_S2
  `define AXI_R_LAYER_M13_S2 `i_axi_AXI_R_LAYER_M13_S2
`endif 

`ifdef i_axi_AXI_R_LAYER_M13_S3
  `define AXI_R_LAYER_M13_S3 `i_axi_AXI_R_LAYER_M13_S3
`endif 

`ifdef i_axi_AXI_R_LAYER_M13_S4
  `define AXI_R_LAYER_M13_S4 `i_axi_AXI_R_LAYER_M13_S4
`endif 

`ifdef i_axi_AXI_R_LAYER_M13_S5
  `define AXI_R_LAYER_M13_S5 `i_axi_AXI_R_LAYER_M13_S5
`endif 

`ifdef i_axi_AXI_R_LAYER_M13_S6
  `define AXI_R_LAYER_M13_S6 `i_axi_AXI_R_LAYER_M13_S6
`endif 

`ifdef i_axi_AXI_R_LAYER_M13_S7
  `define AXI_R_LAYER_M13_S7 `i_axi_AXI_R_LAYER_M13_S7
`endif 

`ifdef i_axi_AXI_R_LAYER_M13_S8
  `define AXI_R_LAYER_M13_S8 `i_axi_AXI_R_LAYER_M13_S8
`endif 

`ifdef i_axi_AXI_R_LAYER_M13_S9
  `define AXI_R_LAYER_M13_S9 `i_axi_AXI_R_LAYER_M13_S9
`endif 

`ifdef i_axi_AXI_R_LAYER_M13_S10
  `define AXI_R_LAYER_M13_S10 `i_axi_AXI_R_LAYER_M13_S10
`endif 

`ifdef i_axi_AXI_R_LAYER_M13_S11
  `define AXI_R_LAYER_M13_S11 `i_axi_AXI_R_LAYER_M13_S11
`endif 

`ifdef i_axi_AXI_R_LAYER_M13_S12
  `define AXI_R_LAYER_M13_S12 `i_axi_AXI_R_LAYER_M13_S12
`endif 

`ifdef i_axi_AXI_R_LAYER_M13_S13
  `define AXI_R_LAYER_M13_S13 `i_axi_AXI_R_LAYER_M13_S13
`endif 

`ifdef i_axi_AXI_R_LAYER_M13_S14
  `define AXI_R_LAYER_M13_S14 `i_axi_AXI_R_LAYER_M13_S14
`endif 

`ifdef i_axi_AXI_R_LAYER_M13_S15
  `define AXI_R_LAYER_M13_S15 `i_axi_AXI_R_LAYER_M13_S15
`endif 

`ifdef i_axi_AXI_R_LAYER_M13_S16
  `define AXI_R_LAYER_M13_S16 `i_axi_AXI_R_LAYER_M13_S16
`endif 

`ifdef i_axi_AXI_B_LAYER_M13_S0
  `define AXI_B_LAYER_M13_S0 `i_axi_AXI_B_LAYER_M13_S0
`endif 

`ifdef i_axi_AXI_B_LAYER_M13_S1
  `define AXI_B_LAYER_M13_S1 `i_axi_AXI_B_LAYER_M13_S1
`endif 

`ifdef i_axi_AXI_B_LAYER_M13_S2
  `define AXI_B_LAYER_M13_S2 `i_axi_AXI_B_LAYER_M13_S2
`endif 

`ifdef i_axi_AXI_B_LAYER_M13_S3
  `define AXI_B_LAYER_M13_S3 `i_axi_AXI_B_LAYER_M13_S3
`endif 

`ifdef i_axi_AXI_B_LAYER_M13_S4
  `define AXI_B_LAYER_M13_S4 `i_axi_AXI_B_LAYER_M13_S4
`endif 

`ifdef i_axi_AXI_B_LAYER_M13_S5
  `define AXI_B_LAYER_M13_S5 `i_axi_AXI_B_LAYER_M13_S5
`endif 

`ifdef i_axi_AXI_B_LAYER_M13_S6
  `define AXI_B_LAYER_M13_S6 `i_axi_AXI_B_LAYER_M13_S6
`endif 

`ifdef i_axi_AXI_B_LAYER_M13_S7
  `define AXI_B_LAYER_M13_S7 `i_axi_AXI_B_LAYER_M13_S7
`endif 

`ifdef i_axi_AXI_B_LAYER_M13_S8
  `define AXI_B_LAYER_M13_S8 `i_axi_AXI_B_LAYER_M13_S8
`endif 

`ifdef i_axi_AXI_B_LAYER_M13_S9
  `define AXI_B_LAYER_M13_S9 `i_axi_AXI_B_LAYER_M13_S9
`endif 

`ifdef i_axi_AXI_B_LAYER_M13_S10
  `define AXI_B_LAYER_M13_S10 `i_axi_AXI_B_LAYER_M13_S10
`endif 

`ifdef i_axi_AXI_B_LAYER_M13_S11
  `define AXI_B_LAYER_M13_S11 `i_axi_AXI_B_LAYER_M13_S11
`endif 

`ifdef i_axi_AXI_B_LAYER_M13_S12
  `define AXI_B_LAYER_M13_S12 `i_axi_AXI_B_LAYER_M13_S12
`endif 

`ifdef i_axi_AXI_B_LAYER_M13_S13
  `define AXI_B_LAYER_M13_S13 `i_axi_AXI_B_LAYER_M13_S13
`endif 

`ifdef i_axi_AXI_B_LAYER_M13_S14
  `define AXI_B_LAYER_M13_S14 `i_axi_AXI_B_LAYER_M13_S14
`endif 

`ifdef i_axi_AXI_B_LAYER_M13_S15
  `define AXI_B_LAYER_M13_S15 `i_axi_AXI_B_LAYER_M13_S15
`endif 

`ifdef i_axi_AXI_B_LAYER_M13_S16
  `define AXI_B_LAYER_M13_S16 `i_axi_AXI_B_LAYER_M13_S16
`endif 

`ifdef i_axi_AXI_R_LAYER_M14_S0
  `define AXI_R_LAYER_M14_S0 `i_axi_AXI_R_LAYER_M14_S0
`endif 

`ifdef i_axi_AXI_R_LAYER_M14_S1
  `define AXI_R_LAYER_M14_S1 `i_axi_AXI_R_LAYER_M14_S1
`endif 

`ifdef i_axi_AXI_R_LAYER_M14_S2
  `define AXI_R_LAYER_M14_S2 `i_axi_AXI_R_LAYER_M14_S2
`endif 

`ifdef i_axi_AXI_R_LAYER_M14_S3
  `define AXI_R_LAYER_M14_S3 `i_axi_AXI_R_LAYER_M14_S3
`endif 

`ifdef i_axi_AXI_R_LAYER_M14_S4
  `define AXI_R_LAYER_M14_S4 `i_axi_AXI_R_LAYER_M14_S4
`endif 

`ifdef i_axi_AXI_R_LAYER_M14_S5
  `define AXI_R_LAYER_M14_S5 `i_axi_AXI_R_LAYER_M14_S5
`endif 

`ifdef i_axi_AXI_R_LAYER_M14_S6
  `define AXI_R_LAYER_M14_S6 `i_axi_AXI_R_LAYER_M14_S6
`endif 

`ifdef i_axi_AXI_R_LAYER_M14_S7
  `define AXI_R_LAYER_M14_S7 `i_axi_AXI_R_LAYER_M14_S7
`endif 

`ifdef i_axi_AXI_R_LAYER_M14_S8
  `define AXI_R_LAYER_M14_S8 `i_axi_AXI_R_LAYER_M14_S8
`endif 

`ifdef i_axi_AXI_R_LAYER_M14_S9
  `define AXI_R_LAYER_M14_S9 `i_axi_AXI_R_LAYER_M14_S9
`endif 

`ifdef i_axi_AXI_R_LAYER_M14_S10
  `define AXI_R_LAYER_M14_S10 `i_axi_AXI_R_LAYER_M14_S10
`endif 

`ifdef i_axi_AXI_R_LAYER_M14_S11
  `define AXI_R_LAYER_M14_S11 `i_axi_AXI_R_LAYER_M14_S11
`endif 

`ifdef i_axi_AXI_R_LAYER_M14_S12
  `define AXI_R_LAYER_M14_S12 `i_axi_AXI_R_LAYER_M14_S12
`endif 

`ifdef i_axi_AXI_R_LAYER_M14_S13
  `define AXI_R_LAYER_M14_S13 `i_axi_AXI_R_LAYER_M14_S13
`endif 

`ifdef i_axi_AXI_R_LAYER_M14_S14
  `define AXI_R_LAYER_M14_S14 `i_axi_AXI_R_LAYER_M14_S14
`endif 

`ifdef i_axi_AXI_R_LAYER_M14_S15
  `define AXI_R_LAYER_M14_S15 `i_axi_AXI_R_LAYER_M14_S15
`endif 

`ifdef i_axi_AXI_R_LAYER_M14_S16
  `define AXI_R_LAYER_M14_S16 `i_axi_AXI_R_LAYER_M14_S16
`endif 

`ifdef i_axi_AXI_B_LAYER_M14_S0
  `define AXI_B_LAYER_M14_S0 `i_axi_AXI_B_LAYER_M14_S0
`endif 

`ifdef i_axi_AXI_B_LAYER_M14_S1
  `define AXI_B_LAYER_M14_S1 `i_axi_AXI_B_LAYER_M14_S1
`endif 

`ifdef i_axi_AXI_B_LAYER_M14_S2
  `define AXI_B_LAYER_M14_S2 `i_axi_AXI_B_LAYER_M14_S2
`endif 

`ifdef i_axi_AXI_B_LAYER_M14_S3
  `define AXI_B_LAYER_M14_S3 `i_axi_AXI_B_LAYER_M14_S3
`endif 

`ifdef i_axi_AXI_B_LAYER_M14_S4
  `define AXI_B_LAYER_M14_S4 `i_axi_AXI_B_LAYER_M14_S4
`endif 

`ifdef i_axi_AXI_B_LAYER_M14_S5
  `define AXI_B_LAYER_M14_S5 `i_axi_AXI_B_LAYER_M14_S5
`endif 

`ifdef i_axi_AXI_B_LAYER_M14_S6
  `define AXI_B_LAYER_M14_S6 `i_axi_AXI_B_LAYER_M14_S6
`endif 

`ifdef i_axi_AXI_B_LAYER_M14_S7
  `define AXI_B_LAYER_M14_S7 `i_axi_AXI_B_LAYER_M14_S7
`endif 

`ifdef i_axi_AXI_B_LAYER_M14_S8
  `define AXI_B_LAYER_M14_S8 `i_axi_AXI_B_LAYER_M14_S8
`endif 

`ifdef i_axi_AXI_B_LAYER_M14_S9
  `define AXI_B_LAYER_M14_S9 `i_axi_AXI_B_LAYER_M14_S9
`endif 

`ifdef i_axi_AXI_B_LAYER_M14_S10
  `define AXI_B_LAYER_M14_S10 `i_axi_AXI_B_LAYER_M14_S10
`endif 

`ifdef i_axi_AXI_B_LAYER_M14_S11
  `define AXI_B_LAYER_M14_S11 `i_axi_AXI_B_LAYER_M14_S11
`endif 

`ifdef i_axi_AXI_B_LAYER_M14_S12
  `define AXI_B_LAYER_M14_S12 `i_axi_AXI_B_LAYER_M14_S12
`endif 

`ifdef i_axi_AXI_B_LAYER_M14_S13
  `define AXI_B_LAYER_M14_S13 `i_axi_AXI_B_LAYER_M14_S13
`endif 

`ifdef i_axi_AXI_B_LAYER_M14_S14
  `define AXI_B_LAYER_M14_S14 `i_axi_AXI_B_LAYER_M14_S14
`endif 

`ifdef i_axi_AXI_B_LAYER_M14_S15
  `define AXI_B_LAYER_M14_S15 `i_axi_AXI_B_LAYER_M14_S15
`endif 

`ifdef i_axi_AXI_B_LAYER_M14_S16
  `define AXI_B_LAYER_M14_S16 `i_axi_AXI_B_LAYER_M14_S16
`endif 

`ifdef i_axi_AXI_R_LAYER_M15_S0
  `define AXI_R_LAYER_M15_S0 `i_axi_AXI_R_LAYER_M15_S0
`endif 

`ifdef i_axi_AXI_R_LAYER_M15_S1
  `define AXI_R_LAYER_M15_S1 `i_axi_AXI_R_LAYER_M15_S1
`endif 

`ifdef i_axi_AXI_R_LAYER_M15_S2
  `define AXI_R_LAYER_M15_S2 `i_axi_AXI_R_LAYER_M15_S2
`endif 

`ifdef i_axi_AXI_R_LAYER_M15_S3
  `define AXI_R_LAYER_M15_S3 `i_axi_AXI_R_LAYER_M15_S3
`endif 

`ifdef i_axi_AXI_R_LAYER_M15_S4
  `define AXI_R_LAYER_M15_S4 `i_axi_AXI_R_LAYER_M15_S4
`endif 

`ifdef i_axi_AXI_R_LAYER_M15_S5
  `define AXI_R_LAYER_M15_S5 `i_axi_AXI_R_LAYER_M15_S5
`endif 

`ifdef i_axi_AXI_R_LAYER_M15_S6
  `define AXI_R_LAYER_M15_S6 `i_axi_AXI_R_LAYER_M15_S6
`endif 

`ifdef i_axi_AXI_R_LAYER_M15_S7
  `define AXI_R_LAYER_M15_S7 `i_axi_AXI_R_LAYER_M15_S7
`endif 

`ifdef i_axi_AXI_R_LAYER_M15_S8
  `define AXI_R_LAYER_M15_S8 `i_axi_AXI_R_LAYER_M15_S8
`endif 

`ifdef i_axi_AXI_R_LAYER_M15_S9
  `define AXI_R_LAYER_M15_S9 `i_axi_AXI_R_LAYER_M15_S9
`endif 

`ifdef i_axi_AXI_R_LAYER_M15_S10
  `define AXI_R_LAYER_M15_S10 `i_axi_AXI_R_LAYER_M15_S10
`endif 

`ifdef i_axi_AXI_R_LAYER_M15_S11
  `define AXI_R_LAYER_M15_S11 `i_axi_AXI_R_LAYER_M15_S11
`endif 

`ifdef i_axi_AXI_R_LAYER_M15_S12
  `define AXI_R_LAYER_M15_S12 `i_axi_AXI_R_LAYER_M15_S12
`endif 

`ifdef i_axi_AXI_R_LAYER_M15_S13
  `define AXI_R_LAYER_M15_S13 `i_axi_AXI_R_LAYER_M15_S13
`endif 

`ifdef i_axi_AXI_R_LAYER_M15_S14
  `define AXI_R_LAYER_M15_S14 `i_axi_AXI_R_LAYER_M15_S14
`endif 

`ifdef i_axi_AXI_R_LAYER_M15_S15
  `define AXI_R_LAYER_M15_S15 `i_axi_AXI_R_LAYER_M15_S15
`endif 

`ifdef i_axi_AXI_R_LAYER_M15_S16
  `define AXI_R_LAYER_M15_S16 `i_axi_AXI_R_LAYER_M15_S16
`endif 

`ifdef i_axi_AXI_B_LAYER_M15_S0
  `define AXI_B_LAYER_M15_S0 `i_axi_AXI_B_LAYER_M15_S0
`endif 

`ifdef i_axi_AXI_B_LAYER_M15_S1
  `define AXI_B_LAYER_M15_S1 `i_axi_AXI_B_LAYER_M15_S1
`endif 

`ifdef i_axi_AXI_B_LAYER_M15_S2
  `define AXI_B_LAYER_M15_S2 `i_axi_AXI_B_LAYER_M15_S2
`endif 

`ifdef i_axi_AXI_B_LAYER_M15_S3
  `define AXI_B_LAYER_M15_S3 `i_axi_AXI_B_LAYER_M15_S3
`endif 

`ifdef i_axi_AXI_B_LAYER_M15_S4
  `define AXI_B_LAYER_M15_S4 `i_axi_AXI_B_LAYER_M15_S4
`endif 

`ifdef i_axi_AXI_B_LAYER_M15_S5
  `define AXI_B_LAYER_M15_S5 `i_axi_AXI_B_LAYER_M15_S5
`endif 

`ifdef i_axi_AXI_B_LAYER_M15_S6
  `define AXI_B_LAYER_M15_S6 `i_axi_AXI_B_LAYER_M15_S6
`endif 

`ifdef i_axi_AXI_B_LAYER_M15_S7
  `define AXI_B_LAYER_M15_S7 `i_axi_AXI_B_LAYER_M15_S7
`endif 

`ifdef i_axi_AXI_B_LAYER_M15_S8
  `define AXI_B_LAYER_M15_S8 `i_axi_AXI_B_LAYER_M15_S8
`endif 

`ifdef i_axi_AXI_B_LAYER_M15_S9
  `define AXI_B_LAYER_M15_S9 `i_axi_AXI_B_LAYER_M15_S9
`endif 

`ifdef i_axi_AXI_B_LAYER_M15_S10
  `define AXI_B_LAYER_M15_S10 `i_axi_AXI_B_LAYER_M15_S10
`endif 

`ifdef i_axi_AXI_B_LAYER_M15_S11
  `define AXI_B_LAYER_M15_S11 `i_axi_AXI_B_LAYER_M15_S11
`endif 

`ifdef i_axi_AXI_B_LAYER_M15_S12
  `define AXI_B_LAYER_M15_S12 `i_axi_AXI_B_LAYER_M15_S12
`endif 

`ifdef i_axi_AXI_B_LAYER_M15_S13
  `define AXI_B_LAYER_M15_S13 `i_axi_AXI_B_LAYER_M15_S13
`endif 

`ifdef i_axi_AXI_B_LAYER_M15_S14
  `define AXI_B_LAYER_M15_S14 `i_axi_AXI_B_LAYER_M15_S14
`endif 

`ifdef i_axi_AXI_B_LAYER_M15_S15
  `define AXI_B_LAYER_M15_S15 `i_axi_AXI_B_LAYER_M15_S15
`endif 

`ifdef i_axi_AXI_B_LAYER_M15_S16
  `define AXI_B_LAYER_M15_S16 `i_axi_AXI_B_LAYER_M15_S16
`endif 

`ifdef i_axi_AXI_R_LAYER_M16_S0
  `define AXI_R_LAYER_M16_S0 `i_axi_AXI_R_LAYER_M16_S0
`endif 

`ifdef i_axi_AXI_R_LAYER_M16_S1
  `define AXI_R_LAYER_M16_S1 `i_axi_AXI_R_LAYER_M16_S1
`endif 

`ifdef i_axi_AXI_R_LAYER_M16_S2
  `define AXI_R_LAYER_M16_S2 `i_axi_AXI_R_LAYER_M16_S2
`endif 

`ifdef i_axi_AXI_R_LAYER_M16_S3
  `define AXI_R_LAYER_M16_S3 `i_axi_AXI_R_LAYER_M16_S3
`endif 

`ifdef i_axi_AXI_R_LAYER_M16_S4
  `define AXI_R_LAYER_M16_S4 `i_axi_AXI_R_LAYER_M16_S4
`endif 

`ifdef i_axi_AXI_R_LAYER_M16_S5
  `define AXI_R_LAYER_M16_S5 `i_axi_AXI_R_LAYER_M16_S5
`endif 

`ifdef i_axi_AXI_R_LAYER_M16_S6
  `define AXI_R_LAYER_M16_S6 `i_axi_AXI_R_LAYER_M16_S6
`endif 

`ifdef i_axi_AXI_R_LAYER_M16_S7
  `define AXI_R_LAYER_M16_S7 `i_axi_AXI_R_LAYER_M16_S7
`endif 

`ifdef i_axi_AXI_R_LAYER_M16_S8
  `define AXI_R_LAYER_M16_S8 `i_axi_AXI_R_LAYER_M16_S8
`endif 

`ifdef i_axi_AXI_R_LAYER_M16_S9
  `define AXI_R_LAYER_M16_S9 `i_axi_AXI_R_LAYER_M16_S9
`endif 

`ifdef i_axi_AXI_R_LAYER_M16_S10
  `define AXI_R_LAYER_M16_S10 `i_axi_AXI_R_LAYER_M16_S10
`endif 

`ifdef i_axi_AXI_R_LAYER_M16_S11
  `define AXI_R_LAYER_M16_S11 `i_axi_AXI_R_LAYER_M16_S11
`endif 

`ifdef i_axi_AXI_R_LAYER_M16_S12
  `define AXI_R_LAYER_M16_S12 `i_axi_AXI_R_LAYER_M16_S12
`endif 

`ifdef i_axi_AXI_R_LAYER_M16_S13
  `define AXI_R_LAYER_M16_S13 `i_axi_AXI_R_LAYER_M16_S13
`endif 

`ifdef i_axi_AXI_R_LAYER_M16_S14
  `define AXI_R_LAYER_M16_S14 `i_axi_AXI_R_LAYER_M16_S14
`endif 

`ifdef i_axi_AXI_R_LAYER_M16_S15
  `define AXI_R_LAYER_M16_S15 `i_axi_AXI_R_LAYER_M16_S15
`endif 

`ifdef i_axi_AXI_R_LAYER_M16_S16
  `define AXI_R_LAYER_M16_S16 `i_axi_AXI_R_LAYER_M16_S16
`endif 

`ifdef i_axi_AXI_B_LAYER_M16_S0
  `define AXI_B_LAYER_M16_S0 `i_axi_AXI_B_LAYER_M16_S0
`endif 

`ifdef i_axi_AXI_B_LAYER_M16_S1
  `define AXI_B_LAYER_M16_S1 `i_axi_AXI_B_LAYER_M16_S1
`endif 

`ifdef i_axi_AXI_B_LAYER_M16_S2
  `define AXI_B_LAYER_M16_S2 `i_axi_AXI_B_LAYER_M16_S2
`endif 

`ifdef i_axi_AXI_B_LAYER_M16_S3
  `define AXI_B_LAYER_M16_S3 `i_axi_AXI_B_LAYER_M16_S3
`endif 

`ifdef i_axi_AXI_B_LAYER_M16_S4
  `define AXI_B_LAYER_M16_S4 `i_axi_AXI_B_LAYER_M16_S4
`endif 

`ifdef i_axi_AXI_B_LAYER_M16_S5
  `define AXI_B_LAYER_M16_S5 `i_axi_AXI_B_LAYER_M16_S5
`endif 

`ifdef i_axi_AXI_B_LAYER_M16_S6
  `define AXI_B_LAYER_M16_S6 `i_axi_AXI_B_LAYER_M16_S6
`endif 

`ifdef i_axi_AXI_B_LAYER_M16_S7
  `define AXI_B_LAYER_M16_S7 `i_axi_AXI_B_LAYER_M16_S7
`endif 

`ifdef i_axi_AXI_B_LAYER_M16_S8
  `define AXI_B_LAYER_M16_S8 `i_axi_AXI_B_LAYER_M16_S8
`endif 

`ifdef i_axi_AXI_B_LAYER_M16_S9
  `define AXI_B_LAYER_M16_S9 `i_axi_AXI_B_LAYER_M16_S9
`endif 

`ifdef i_axi_AXI_B_LAYER_M16_S10
  `define AXI_B_LAYER_M16_S10 `i_axi_AXI_B_LAYER_M16_S10
`endif 

`ifdef i_axi_AXI_B_LAYER_M16_S11
  `define AXI_B_LAYER_M16_S11 `i_axi_AXI_B_LAYER_M16_S11
`endif 

`ifdef i_axi_AXI_B_LAYER_M16_S12
  `define AXI_B_LAYER_M16_S12 `i_axi_AXI_B_LAYER_M16_S12
`endif 

`ifdef i_axi_AXI_B_LAYER_M16_S13
  `define AXI_B_LAYER_M16_S13 `i_axi_AXI_B_LAYER_M16_S13
`endif 

`ifdef i_axi_AXI_B_LAYER_M16_S14
  `define AXI_B_LAYER_M16_S14 `i_axi_AXI_B_LAYER_M16_S14
`endif 

`ifdef i_axi_AXI_B_LAYER_M16_S15
  `define AXI_B_LAYER_M16_S15 `i_axi_AXI_B_LAYER_M16_S15
`endif 

`ifdef i_axi_AXI_B_LAYER_M16_S16
  `define AXI_B_LAYER_M16_S16 `i_axi_AXI_B_LAYER_M16_S16
`endif 

`ifdef i_axi_AXI_AR_HAS_SHARED_LAYER
  `define AXI_AR_HAS_SHARED_LAYER `i_axi_AXI_AR_HAS_SHARED_LAYER
`endif 

`ifdef i_axi_AXI_AR_SHARED_LAYER
  `define AXI_AR_SHARED_LAYER `i_axi_AXI_AR_SHARED_LAYER
`endif 

`ifdef i_axi_AXI_AW_HAS_SHARED_LAYER
  `define AXI_AW_HAS_SHARED_LAYER `i_axi_AXI_AW_HAS_SHARED_LAYER
`endif 

`ifdef i_axi_AXI_AW_SHARED_LAYER
  `define AXI_AW_SHARED_LAYER `i_axi_AXI_AW_SHARED_LAYER
`endif 

`ifdef i_axi_AXI_W_HAS_SHARED_LAYER
  `define AXI_W_HAS_SHARED_LAYER `i_axi_AXI_W_HAS_SHARED_LAYER
`endif 

`ifdef i_axi_AXI_W_SHARED_LAYER
  `define AXI_W_SHARED_LAYER `i_axi_AXI_W_SHARED_LAYER
`endif 

`ifdef i_axi_AXI_R_HAS_SHARED_LAYER
  `define AXI_R_HAS_SHARED_LAYER `i_axi_AXI_R_HAS_SHARED_LAYER
`endif 

`ifdef i_axi_AXI_R_SHARED_LAYER
  `define AXI_R_SHARED_LAYER `i_axi_AXI_R_SHARED_LAYER
`endif 

`ifdef i_axi_AXI_B_HAS_SHARED_LAYER
  `define AXI_B_HAS_SHARED_LAYER `i_axi_AXI_B_HAS_SHARED_LAYER
`endif 

`ifdef i_axi_AXI_B_SHARED_LAYER
  `define AXI_B_SHARED_LAYER `i_axi_AXI_B_SHARED_LAYER
`endif 

`ifdef i_axi_AXI_AR_SHARED_LAYER_NM
  `define AXI_AR_SHARED_LAYER_NM `i_axi_AXI_AR_SHARED_LAYER_NM
`endif 

`ifdef i_axi_AXI_LOG2_AR_SHARED_LAYER_NM
  `define AXI_LOG2_AR_SHARED_LAYER_NM `i_axi_AXI_LOG2_AR_SHARED_LAYER_NM
`endif 

`ifdef i_axi_AXI_LOG2_AR_SHARED_LAYER_NMP1
  `define AXI_LOG2_AR_SHARED_LAYER_NMP1 `i_axi_AXI_LOG2_AR_SHARED_LAYER_NMP1
`endif 

`ifdef i_axi_AXI_AR_SHARED_LAYER_NS
  `define AXI_AR_SHARED_LAYER_NS `i_axi_AXI_AR_SHARED_LAYER_NS
`endif 

`ifdef i_axi_AXI_AR_SHARED_LAYER_NS_R0
  `define AXI_AR_SHARED_LAYER_NS_R0 `i_axi_AXI_AR_SHARED_LAYER_NS_R0
`endif 

`ifdef i_axi_AXI_LOG2_AR_SHARED_LAYER_NS
  `define AXI_LOG2_AR_SHARED_LAYER_NS `i_axi_AXI_LOG2_AR_SHARED_LAYER_NS
`endif 

`ifdef i_axi_AXI_LOG2_AR_SHARED_LAYER_NSP1
  `define AXI_LOG2_AR_SHARED_LAYER_NSP1 `i_axi_AXI_LOG2_AR_SHARED_LAYER_NSP1
`endif 

`ifdef i_axi_AXI_AW_SHARED_LAYER_NM
  `define AXI_AW_SHARED_LAYER_NM `i_axi_AXI_AW_SHARED_LAYER_NM
`endif 

`ifdef i_axi_AXI_LOG2_AW_SHARED_LAYER_NM
  `define AXI_LOG2_AW_SHARED_LAYER_NM `i_axi_AXI_LOG2_AW_SHARED_LAYER_NM
`endif 

`ifdef i_axi_AXI_LOG2_AW_SHARED_LAYER_NMP1
  `define AXI_LOG2_AW_SHARED_LAYER_NMP1 `i_axi_AXI_LOG2_AW_SHARED_LAYER_NMP1
`endif 

`ifdef i_axi_AXI_AW_SHARED_LAYER_NS
  `define AXI_AW_SHARED_LAYER_NS `i_axi_AXI_AW_SHARED_LAYER_NS
`endif 

`ifdef i_axi_AXI_AW_SHARED_LAYER_NS_R0
  `define AXI_AW_SHARED_LAYER_NS_R0 `i_axi_AXI_AW_SHARED_LAYER_NS_R0
`endif 

`ifdef i_axi_AXI_LOG2_AW_SHARED_LAYER_NS
  `define AXI_LOG2_AW_SHARED_LAYER_NS `i_axi_AXI_LOG2_AW_SHARED_LAYER_NS
`endif 

`ifdef i_axi_AXI_LOG2_AW_SHARED_LAYER_NSP1
  `define AXI_LOG2_AW_SHARED_LAYER_NSP1 `i_axi_AXI_LOG2_AW_SHARED_LAYER_NSP1
`endif 

`ifdef i_axi_AXI_W_SHARED_LAYER_NM
  `define AXI_W_SHARED_LAYER_NM `i_axi_AXI_W_SHARED_LAYER_NM
`endif 

`ifdef i_axi_AXI_LOG2_W_SHARED_LAYER_NM
  `define AXI_LOG2_W_SHARED_LAYER_NM `i_axi_AXI_LOG2_W_SHARED_LAYER_NM
`endif 

`ifdef i_axi_AXI_LOG2_W_SHARED_LAYER_NMP1
  `define AXI_LOG2_W_SHARED_LAYER_NMP1 `i_axi_AXI_LOG2_W_SHARED_LAYER_NMP1
`endif 

`ifdef i_axi_AXI_W_SHARED_LAYER_NS
  `define AXI_W_SHARED_LAYER_NS `i_axi_AXI_W_SHARED_LAYER_NS
`endif 

`ifdef i_axi_AXI_W_SHARED_LAYER_NS_R0
  `define AXI_W_SHARED_LAYER_NS_R0 `i_axi_AXI_W_SHARED_LAYER_NS_R0
`endif 

`ifdef i_axi_AXI_LOG2_W_SHARED_LAYER_NS
  `define AXI_LOG2_W_SHARED_LAYER_NS `i_axi_AXI_LOG2_W_SHARED_LAYER_NS
`endif 

`ifdef i_axi_AXI_LOG2_W_SHARED_LAYER_NSP1
  `define AXI_LOG2_W_SHARED_LAYER_NSP1 `i_axi_AXI_LOG2_W_SHARED_LAYER_NSP1
`endif 

`ifdef i_axi_AXI_R_SHARED_LAYER_NM
  `define AXI_R_SHARED_LAYER_NM `i_axi_AXI_R_SHARED_LAYER_NM
`endif 

`ifdef i_axi_AXI_R_SHARED_LAYER_NM_R0
  `define AXI_R_SHARED_LAYER_NM_R0 `i_axi_AXI_R_SHARED_LAYER_NM_R0
`endif 

`ifdef i_axi_AXI_LOG2_R_SHARED_LAYER_NM
  `define AXI_LOG2_R_SHARED_LAYER_NM `i_axi_AXI_LOG2_R_SHARED_LAYER_NM
`endif 

`ifdef i_axi_AXI_LOG2_R_SHARED_LAYER_NMP1
  `define AXI_LOG2_R_SHARED_LAYER_NMP1 `i_axi_AXI_LOG2_R_SHARED_LAYER_NMP1
`endif 

`ifdef i_axi_AXI_R_SHARED_LAYER_NS
  `define AXI_R_SHARED_LAYER_NS `i_axi_AXI_R_SHARED_LAYER_NS
`endif 

`ifdef i_axi_AXI_LOG2_R_SHARED_LAYER_NS
  `define AXI_LOG2_R_SHARED_LAYER_NS `i_axi_AXI_LOG2_R_SHARED_LAYER_NS
`endif 

`ifdef i_axi_AXI_LOG2_R_SHARED_LAYER_NSP1
  `define AXI_LOG2_R_SHARED_LAYER_NSP1 `i_axi_AXI_LOG2_R_SHARED_LAYER_NSP1
`endif 

`ifdef i_axi_AXI_B_SHARED_LAYER_NM
  `define AXI_B_SHARED_LAYER_NM `i_axi_AXI_B_SHARED_LAYER_NM
`endif 

`ifdef i_axi_AXI_B_SHARED_LAYER_NM_R0
  `define AXI_B_SHARED_LAYER_NM_R0 `i_axi_AXI_B_SHARED_LAYER_NM_R0
`endif 

`ifdef i_axi_AXI_LOG2_B_SHARED_LAYER_NM
  `define AXI_LOG2_B_SHARED_LAYER_NM `i_axi_AXI_LOG2_B_SHARED_LAYER_NM
`endif 

`ifdef i_axi_AXI_LOG2_B_SHARED_LAYER_NMP1
  `define AXI_LOG2_B_SHARED_LAYER_NMP1 `i_axi_AXI_LOG2_B_SHARED_LAYER_NMP1
`endif 

`ifdef i_axi_AXI_B_SHARED_LAYER_NS
  `define AXI_B_SHARED_LAYER_NS `i_axi_AXI_B_SHARED_LAYER_NS
`endif 

`ifdef i_axi_AXI_LOG2_B_SHARED_LAYER_NS
  `define AXI_LOG2_B_SHARED_LAYER_NS `i_axi_AXI_LOG2_B_SHARED_LAYER_NS
`endif 

`ifdef i_axi_AXI_LOG2_B_SHARED_LAYER_NSP1
  `define AXI_LOG2_B_SHARED_LAYER_NSP1 `i_axi_AXI_LOG2_B_SHARED_LAYER_NSP1
`endif 

`ifdef i_axi_AXI_AR_S0_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AR_S0_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AR_S0_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AR_S0_HAS_SHRD_DDCTD_LNK
  `define AXI_AR_S0_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AR_S0_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AR_S0_NMV
  `define AXI_AR_S0_NMV `i_axi_AXI_AR_S0_NMV
`endif 

`ifdef i_axi_AXI_AR_S0_NMV_LOG2
  `define AXI_AR_S0_NMV_LOG2 `i_axi_AXI_AR_S0_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AR_S0_NMV_P1_LOG2
  `define AXI_AR_S0_NMV_P1_LOG2 `i_axi_AXI_AR_S0_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AW_S0_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AW_S0_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AW_S0_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AW_S0_HAS_SHRD_DDCTD_LNK
  `define AXI_AW_S0_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AW_S0_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AW_S0_NMV
  `define AXI_AW_S0_NMV `i_axi_AXI_AW_S0_NMV
`endif 

`ifdef i_axi_AXI_AW_S0_NMV_LOG2
  `define AXI_AW_S0_NMV_LOG2 `i_axi_AXI_AW_S0_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AW_S0_NMV_P1_LOG2
  `define AXI_AW_S0_NMV_P1_LOG2 `i_axi_AXI_AW_S0_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_W_S0_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_W_S0_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_W_S0_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_W_S0_HAS_SHRD_DDCTD_LNK
  `define AXI_W_S0_HAS_SHRD_DDCTD_LNK `i_axi_AXI_W_S0_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_W_S0_NMV
  `define AXI_W_S0_NMV `i_axi_AXI_W_S0_NMV
`endif 

`ifdef i_axi_AXI_W_S0_NMV_LOG2
  `define AXI_W_S0_NMV_LOG2 `i_axi_AXI_W_S0_NMV_LOG2
`endif 

`ifdef i_axi_AXI_W_S0_NMV_P1_LOG2
  `define AXI_W_S0_NMV_P1_LOG2 `i_axi_AXI_W_S0_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AR_S1_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AR_S1_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AR_S1_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AR_S1_HAS_SHRD_DDCTD_LNK
  `define AXI_AR_S1_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AR_S1_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AR_S1_NMV
  `define AXI_AR_S1_NMV `i_axi_AXI_AR_S1_NMV
`endif 

`ifdef i_axi_AXI_AR_S1_NMV_LOG2
  `define AXI_AR_S1_NMV_LOG2 `i_axi_AXI_AR_S1_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AR_S1_NMV_P1_LOG2
  `define AXI_AR_S1_NMV_P1_LOG2 `i_axi_AXI_AR_S1_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AW_S1_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AW_S1_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AW_S1_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AW_S1_HAS_SHRD_DDCTD_LNK
  `define AXI_AW_S1_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AW_S1_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AW_S1_NMV
  `define AXI_AW_S1_NMV `i_axi_AXI_AW_S1_NMV
`endif 

`ifdef i_axi_AXI_AW_S1_NMV_LOG2
  `define AXI_AW_S1_NMV_LOG2 `i_axi_AXI_AW_S1_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AW_S1_NMV_P1_LOG2
  `define AXI_AW_S1_NMV_P1_LOG2 `i_axi_AXI_AW_S1_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_W_S1_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_W_S1_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_W_S1_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_W_S1_HAS_SHRD_DDCTD_LNK
  `define AXI_W_S1_HAS_SHRD_DDCTD_LNK `i_axi_AXI_W_S1_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_W_S1_NMV
  `define AXI_W_S1_NMV `i_axi_AXI_W_S1_NMV
`endif 

`ifdef i_axi_AXI_W_S1_NMV_LOG2
  `define AXI_W_S1_NMV_LOG2 `i_axi_AXI_W_S1_NMV_LOG2
`endif 

`ifdef i_axi_AXI_W_S1_NMV_P1_LOG2
  `define AXI_W_S1_NMV_P1_LOG2 `i_axi_AXI_W_S1_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AR_S2_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AR_S2_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AR_S2_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AR_S2_HAS_SHRD_DDCTD_LNK
  `define AXI_AR_S2_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AR_S2_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AR_S2_NMV
  `define AXI_AR_S2_NMV `i_axi_AXI_AR_S2_NMV
`endif 

`ifdef i_axi_AXI_AR_S2_NMV_LOG2
  `define AXI_AR_S2_NMV_LOG2 `i_axi_AXI_AR_S2_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AR_S2_NMV_P1_LOG2
  `define AXI_AR_S2_NMV_P1_LOG2 `i_axi_AXI_AR_S2_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AW_S2_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AW_S2_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AW_S2_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AW_S2_HAS_SHRD_DDCTD_LNK
  `define AXI_AW_S2_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AW_S2_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AW_S2_NMV
  `define AXI_AW_S2_NMV `i_axi_AXI_AW_S2_NMV
`endif 

`ifdef i_axi_AXI_AW_S2_NMV_LOG2
  `define AXI_AW_S2_NMV_LOG2 `i_axi_AXI_AW_S2_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AW_S2_NMV_P1_LOG2
  `define AXI_AW_S2_NMV_P1_LOG2 `i_axi_AXI_AW_S2_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_W_S2_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_W_S2_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_W_S2_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_W_S2_HAS_SHRD_DDCTD_LNK
  `define AXI_W_S2_HAS_SHRD_DDCTD_LNK `i_axi_AXI_W_S2_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_W_S2_NMV
  `define AXI_W_S2_NMV `i_axi_AXI_W_S2_NMV
`endif 

`ifdef i_axi_AXI_W_S2_NMV_LOG2
  `define AXI_W_S2_NMV_LOG2 `i_axi_AXI_W_S2_NMV_LOG2
`endif 

`ifdef i_axi_AXI_W_S2_NMV_P1_LOG2
  `define AXI_W_S2_NMV_P1_LOG2 `i_axi_AXI_W_S2_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AR_S3_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AR_S3_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AR_S3_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AR_S3_HAS_SHRD_DDCTD_LNK
  `define AXI_AR_S3_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AR_S3_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AR_S3_NMV
  `define AXI_AR_S3_NMV `i_axi_AXI_AR_S3_NMV
`endif 

`ifdef i_axi_AXI_AR_S3_NMV_LOG2
  `define AXI_AR_S3_NMV_LOG2 `i_axi_AXI_AR_S3_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AR_S3_NMV_P1_LOG2
  `define AXI_AR_S3_NMV_P1_LOG2 `i_axi_AXI_AR_S3_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AW_S3_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AW_S3_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AW_S3_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AW_S3_HAS_SHRD_DDCTD_LNK
  `define AXI_AW_S3_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AW_S3_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AW_S3_NMV
  `define AXI_AW_S3_NMV `i_axi_AXI_AW_S3_NMV
`endif 

`ifdef i_axi_AXI_AW_S3_NMV_LOG2
  `define AXI_AW_S3_NMV_LOG2 `i_axi_AXI_AW_S3_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AW_S3_NMV_P1_LOG2
  `define AXI_AW_S3_NMV_P1_LOG2 `i_axi_AXI_AW_S3_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_W_S3_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_W_S3_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_W_S3_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_W_S3_HAS_SHRD_DDCTD_LNK
  `define AXI_W_S3_HAS_SHRD_DDCTD_LNK `i_axi_AXI_W_S3_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_W_S3_NMV
  `define AXI_W_S3_NMV `i_axi_AXI_W_S3_NMV
`endif 

`ifdef i_axi_AXI_W_S3_NMV_LOG2
  `define AXI_W_S3_NMV_LOG2 `i_axi_AXI_W_S3_NMV_LOG2
`endif 

`ifdef i_axi_AXI_W_S3_NMV_P1_LOG2
  `define AXI_W_S3_NMV_P1_LOG2 `i_axi_AXI_W_S3_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AR_S4_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AR_S4_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AR_S4_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AR_S4_HAS_SHRD_DDCTD_LNK
  `define AXI_AR_S4_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AR_S4_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AR_S4_NMV
  `define AXI_AR_S4_NMV `i_axi_AXI_AR_S4_NMV
`endif 

`ifdef i_axi_AXI_AR_S4_NMV_LOG2
  `define AXI_AR_S4_NMV_LOG2 `i_axi_AXI_AR_S4_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AR_S4_NMV_P1_LOG2
  `define AXI_AR_S4_NMV_P1_LOG2 `i_axi_AXI_AR_S4_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AW_S4_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AW_S4_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AW_S4_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AW_S4_HAS_SHRD_DDCTD_LNK
  `define AXI_AW_S4_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AW_S4_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AW_S4_NMV
  `define AXI_AW_S4_NMV `i_axi_AXI_AW_S4_NMV
`endif 

`ifdef i_axi_AXI_AW_S4_NMV_LOG2
  `define AXI_AW_S4_NMV_LOG2 `i_axi_AXI_AW_S4_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AW_S4_NMV_P1_LOG2
  `define AXI_AW_S4_NMV_P1_LOG2 `i_axi_AXI_AW_S4_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_W_S4_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_W_S4_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_W_S4_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_W_S4_HAS_SHRD_DDCTD_LNK
  `define AXI_W_S4_HAS_SHRD_DDCTD_LNK `i_axi_AXI_W_S4_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_W_S4_NMV
  `define AXI_W_S4_NMV `i_axi_AXI_W_S4_NMV
`endif 

`ifdef i_axi_AXI_W_S4_NMV_LOG2
  `define AXI_W_S4_NMV_LOG2 `i_axi_AXI_W_S4_NMV_LOG2
`endif 

`ifdef i_axi_AXI_W_S4_NMV_P1_LOG2
  `define AXI_W_S4_NMV_P1_LOG2 `i_axi_AXI_W_S4_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AR_S5_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AR_S5_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AR_S5_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AR_S5_HAS_SHRD_DDCTD_LNK
  `define AXI_AR_S5_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AR_S5_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AR_S5_NMV
  `define AXI_AR_S5_NMV `i_axi_AXI_AR_S5_NMV
`endif 

`ifdef i_axi_AXI_AR_S5_NMV_LOG2
  `define AXI_AR_S5_NMV_LOG2 `i_axi_AXI_AR_S5_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AR_S5_NMV_P1_LOG2
  `define AXI_AR_S5_NMV_P1_LOG2 `i_axi_AXI_AR_S5_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AW_S5_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AW_S5_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AW_S5_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AW_S5_HAS_SHRD_DDCTD_LNK
  `define AXI_AW_S5_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AW_S5_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AW_S5_NMV
  `define AXI_AW_S5_NMV `i_axi_AXI_AW_S5_NMV
`endif 

`ifdef i_axi_AXI_AW_S5_NMV_LOG2
  `define AXI_AW_S5_NMV_LOG2 `i_axi_AXI_AW_S5_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AW_S5_NMV_P1_LOG2
  `define AXI_AW_S5_NMV_P1_LOG2 `i_axi_AXI_AW_S5_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_W_S5_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_W_S5_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_W_S5_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_W_S5_HAS_SHRD_DDCTD_LNK
  `define AXI_W_S5_HAS_SHRD_DDCTD_LNK `i_axi_AXI_W_S5_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_W_S5_NMV
  `define AXI_W_S5_NMV `i_axi_AXI_W_S5_NMV
`endif 

`ifdef i_axi_AXI_W_S5_NMV_LOG2
  `define AXI_W_S5_NMV_LOG2 `i_axi_AXI_W_S5_NMV_LOG2
`endif 

`ifdef i_axi_AXI_W_S5_NMV_P1_LOG2
  `define AXI_W_S5_NMV_P1_LOG2 `i_axi_AXI_W_S5_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AR_S6_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AR_S6_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AR_S6_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AR_S6_HAS_SHRD_DDCTD_LNK
  `define AXI_AR_S6_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AR_S6_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AR_S6_NMV
  `define AXI_AR_S6_NMV `i_axi_AXI_AR_S6_NMV
`endif 

`ifdef i_axi_AXI_AR_S6_NMV_LOG2
  `define AXI_AR_S6_NMV_LOG2 `i_axi_AXI_AR_S6_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AR_S6_NMV_P1_LOG2
  `define AXI_AR_S6_NMV_P1_LOG2 `i_axi_AXI_AR_S6_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AW_S6_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AW_S6_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AW_S6_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AW_S6_HAS_SHRD_DDCTD_LNK
  `define AXI_AW_S6_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AW_S6_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AW_S6_NMV
  `define AXI_AW_S6_NMV `i_axi_AXI_AW_S6_NMV
`endif 

`ifdef i_axi_AXI_AW_S6_NMV_LOG2
  `define AXI_AW_S6_NMV_LOG2 `i_axi_AXI_AW_S6_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AW_S6_NMV_P1_LOG2
  `define AXI_AW_S6_NMV_P1_LOG2 `i_axi_AXI_AW_S6_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_W_S6_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_W_S6_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_W_S6_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_W_S6_HAS_SHRD_DDCTD_LNK
  `define AXI_W_S6_HAS_SHRD_DDCTD_LNK `i_axi_AXI_W_S6_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_W_S6_NMV
  `define AXI_W_S6_NMV `i_axi_AXI_W_S6_NMV
`endif 

`ifdef i_axi_AXI_W_S6_NMV_LOG2
  `define AXI_W_S6_NMV_LOG2 `i_axi_AXI_W_S6_NMV_LOG2
`endif 

`ifdef i_axi_AXI_W_S6_NMV_P1_LOG2
  `define AXI_W_S6_NMV_P1_LOG2 `i_axi_AXI_W_S6_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AR_S7_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AR_S7_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AR_S7_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AR_S7_HAS_SHRD_DDCTD_LNK
  `define AXI_AR_S7_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AR_S7_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AR_S7_NMV
  `define AXI_AR_S7_NMV `i_axi_AXI_AR_S7_NMV
`endif 

`ifdef i_axi_AXI_AR_S7_NMV_LOG2
  `define AXI_AR_S7_NMV_LOG2 `i_axi_AXI_AR_S7_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AR_S7_NMV_P1_LOG2
  `define AXI_AR_S7_NMV_P1_LOG2 `i_axi_AXI_AR_S7_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AW_S7_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AW_S7_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AW_S7_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AW_S7_HAS_SHRD_DDCTD_LNK
  `define AXI_AW_S7_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AW_S7_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AW_S7_NMV
  `define AXI_AW_S7_NMV `i_axi_AXI_AW_S7_NMV
`endif 

`ifdef i_axi_AXI_AW_S7_NMV_LOG2
  `define AXI_AW_S7_NMV_LOG2 `i_axi_AXI_AW_S7_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AW_S7_NMV_P1_LOG2
  `define AXI_AW_S7_NMV_P1_LOG2 `i_axi_AXI_AW_S7_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_W_S7_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_W_S7_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_W_S7_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_W_S7_HAS_SHRD_DDCTD_LNK
  `define AXI_W_S7_HAS_SHRD_DDCTD_LNK `i_axi_AXI_W_S7_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_W_S7_NMV
  `define AXI_W_S7_NMV `i_axi_AXI_W_S7_NMV
`endif 

`ifdef i_axi_AXI_W_S7_NMV_LOG2
  `define AXI_W_S7_NMV_LOG2 `i_axi_AXI_W_S7_NMV_LOG2
`endif 

`ifdef i_axi_AXI_W_S7_NMV_P1_LOG2
  `define AXI_W_S7_NMV_P1_LOG2 `i_axi_AXI_W_S7_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AR_S8_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AR_S8_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AR_S8_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AR_S8_HAS_SHRD_DDCTD_LNK
  `define AXI_AR_S8_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AR_S8_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AR_S8_NMV
  `define AXI_AR_S8_NMV `i_axi_AXI_AR_S8_NMV
`endif 

`ifdef i_axi_AXI_AR_S8_NMV_LOG2
  `define AXI_AR_S8_NMV_LOG2 `i_axi_AXI_AR_S8_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AR_S8_NMV_P1_LOG2
  `define AXI_AR_S8_NMV_P1_LOG2 `i_axi_AXI_AR_S8_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AW_S8_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AW_S8_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AW_S8_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AW_S8_HAS_SHRD_DDCTD_LNK
  `define AXI_AW_S8_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AW_S8_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AW_S8_NMV
  `define AXI_AW_S8_NMV `i_axi_AXI_AW_S8_NMV
`endif 

`ifdef i_axi_AXI_AW_S8_NMV_LOG2
  `define AXI_AW_S8_NMV_LOG2 `i_axi_AXI_AW_S8_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AW_S8_NMV_P1_LOG2
  `define AXI_AW_S8_NMV_P1_LOG2 `i_axi_AXI_AW_S8_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_W_S8_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_W_S8_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_W_S8_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_W_S8_HAS_SHRD_DDCTD_LNK
  `define AXI_W_S8_HAS_SHRD_DDCTD_LNK `i_axi_AXI_W_S8_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_W_S8_NMV
  `define AXI_W_S8_NMV `i_axi_AXI_W_S8_NMV
`endif 

`ifdef i_axi_AXI_W_S8_NMV_LOG2
  `define AXI_W_S8_NMV_LOG2 `i_axi_AXI_W_S8_NMV_LOG2
`endif 

`ifdef i_axi_AXI_W_S8_NMV_P1_LOG2
  `define AXI_W_S8_NMV_P1_LOG2 `i_axi_AXI_W_S8_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AR_S9_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AR_S9_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AR_S9_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AR_S9_HAS_SHRD_DDCTD_LNK
  `define AXI_AR_S9_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AR_S9_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AR_S9_NMV
  `define AXI_AR_S9_NMV `i_axi_AXI_AR_S9_NMV
`endif 

`ifdef i_axi_AXI_AR_S9_NMV_LOG2
  `define AXI_AR_S9_NMV_LOG2 `i_axi_AXI_AR_S9_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AR_S9_NMV_P1_LOG2
  `define AXI_AR_S9_NMV_P1_LOG2 `i_axi_AXI_AR_S9_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AW_S9_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AW_S9_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AW_S9_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AW_S9_HAS_SHRD_DDCTD_LNK
  `define AXI_AW_S9_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AW_S9_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AW_S9_NMV
  `define AXI_AW_S9_NMV `i_axi_AXI_AW_S9_NMV
`endif 

`ifdef i_axi_AXI_AW_S9_NMV_LOG2
  `define AXI_AW_S9_NMV_LOG2 `i_axi_AXI_AW_S9_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AW_S9_NMV_P1_LOG2
  `define AXI_AW_S9_NMV_P1_LOG2 `i_axi_AXI_AW_S9_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_W_S9_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_W_S9_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_W_S9_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_W_S9_HAS_SHRD_DDCTD_LNK
  `define AXI_W_S9_HAS_SHRD_DDCTD_LNK `i_axi_AXI_W_S9_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_W_S9_NMV
  `define AXI_W_S9_NMV `i_axi_AXI_W_S9_NMV
`endif 

`ifdef i_axi_AXI_W_S9_NMV_LOG2
  `define AXI_W_S9_NMV_LOG2 `i_axi_AXI_W_S9_NMV_LOG2
`endif 

`ifdef i_axi_AXI_W_S9_NMV_P1_LOG2
  `define AXI_W_S9_NMV_P1_LOG2 `i_axi_AXI_W_S9_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AR_S10_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AR_S10_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AR_S10_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AR_S10_HAS_SHRD_DDCTD_LNK
  `define AXI_AR_S10_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AR_S10_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AR_S10_NMV
  `define AXI_AR_S10_NMV `i_axi_AXI_AR_S10_NMV
`endif 

`ifdef i_axi_AXI_AR_S10_NMV_LOG2
  `define AXI_AR_S10_NMV_LOG2 `i_axi_AXI_AR_S10_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AR_S10_NMV_P1_LOG2
  `define AXI_AR_S10_NMV_P1_LOG2 `i_axi_AXI_AR_S10_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AW_S10_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AW_S10_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AW_S10_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AW_S10_HAS_SHRD_DDCTD_LNK
  `define AXI_AW_S10_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AW_S10_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AW_S10_NMV
  `define AXI_AW_S10_NMV `i_axi_AXI_AW_S10_NMV
`endif 

`ifdef i_axi_AXI_AW_S10_NMV_LOG2
  `define AXI_AW_S10_NMV_LOG2 `i_axi_AXI_AW_S10_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AW_S10_NMV_P1_LOG2
  `define AXI_AW_S10_NMV_P1_LOG2 `i_axi_AXI_AW_S10_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_W_S10_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_W_S10_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_W_S10_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_W_S10_HAS_SHRD_DDCTD_LNK
  `define AXI_W_S10_HAS_SHRD_DDCTD_LNK `i_axi_AXI_W_S10_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_W_S10_NMV
  `define AXI_W_S10_NMV `i_axi_AXI_W_S10_NMV
`endif 

`ifdef i_axi_AXI_W_S10_NMV_LOG2
  `define AXI_W_S10_NMV_LOG2 `i_axi_AXI_W_S10_NMV_LOG2
`endif 

`ifdef i_axi_AXI_W_S10_NMV_P1_LOG2
  `define AXI_W_S10_NMV_P1_LOG2 `i_axi_AXI_W_S10_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AR_S11_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AR_S11_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AR_S11_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AR_S11_HAS_SHRD_DDCTD_LNK
  `define AXI_AR_S11_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AR_S11_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AR_S11_NMV
  `define AXI_AR_S11_NMV `i_axi_AXI_AR_S11_NMV
`endif 

`ifdef i_axi_AXI_AR_S11_NMV_LOG2
  `define AXI_AR_S11_NMV_LOG2 `i_axi_AXI_AR_S11_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AR_S11_NMV_P1_LOG2
  `define AXI_AR_S11_NMV_P1_LOG2 `i_axi_AXI_AR_S11_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AW_S11_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AW_S11_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AW_S11_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AW_S11_HAS_SHRD_DDCTD_LNK
  `define AXI_AW_S11_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AW_S11_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AW_S11_NMV
  `define AXI_AW_S11_NMV `i_axi_AXI_AW_S11_NMV
`endif 

`ifdef i_axi_AXI_AW_S11_NMV_LOG2
  `define AXI_AW_S11_NMV_LOG2 `i_axi_AXI_AW_S11_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AW_S11_NMV_P1_LOG2
  `define AXI_AW_S11_NMV_P1_LOG2 `i_axi_AXI_AW_S11_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_W_S11_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_W_S11_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_W_S11_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_W_S11_HAS_SHRD_DDCTD_LNK
  `define AXI_W_S11_HAS_SHRD_DDCTD_LNK `i_axi_AXI_W_S11_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_W_S11_NMV
  `define AXI_W_S11_NMV `i_axi_AXI_W_S11_NMV
`endif 

`ifdef i_axi_AXI_W_S11_NMV_LOG2
  `define AXI_W_S11_NMV_LOG2 `i_axi_AXI_W_S11_NMV_LOG2
`endif 

`ifdef i_axi_AXI_W_S11_NMV_P1_LOG2
  `define AXI_W_S11_NMV_P1_LOG2 `i_axi_AXI_W_S11_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AR_S12_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AR_S12_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AR_S12_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AR_S12_HAS_SHRD_DDCTD_LNK
  `define AXI_AR_S12_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AR_S12_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AR_S12_NMV
  `define AXI_AR_S12_NMV `i_axi_AXI_AR_S12_NMV
`endif 

`ifdef i_axi_AXI_AR_S12_NMV_LOG2
  `define AXI_AR_S12_NMV_LOG2 `i_axi_AXI_AR_S12_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AR_S12_NMV_P1_LOG2
  `define AXI_AR_S12_NMV_P1_LOG2 `i_axi_AXI_AR_S12_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AW_S12_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AW_S12_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AW_S12_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AW_S12_HAS_SHRD_DDCTD_LNK
  `define AXI_AW_S12_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AW_S12_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AW_S12_NMV
  `define AXI_AW_S12_NMV `i_axi_AXI_AW_S12_NMV
`endif 

`ifdef i_axi_AXI_AW_S12_NMV_LOG2
  `define AXI_AW_S12_NMV_LOG2 `i_axi_AXI_AW_S12_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AW_S12_NMV_P1_LOG2
  `define AXI_AW_S12_NMV_P1_LOG2 `i_axi_AXI_AW_S12_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_W_S12_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_W_S12_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_W_S12_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_W_S12_HAS_SHRD_DDCTD_LNK
  `define AXI_W_S12_HAS_SHRD_DDCTD_LNK `i_axi_AXI_W_S12_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_W_S12_NMV
  `define AXI_W_S12_NMV `i_axi_AXI_W_S12_NMV
`endif 

`ifdef i_axi_AXI_W_S12_NMV_LOG2
  `define AXI_W_S12_NMV_LOG2 `i_axi_AXI_W_S12_NMV_LOG2
`endif 

`ifdef i_axi_AXI_W_S12_NMV_P1_LOG2
  `define AXI_W_S12_NMV_P1_LOG2 `i_axi_AXI_W_S12_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AR_S13_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AR_S13_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AR_S13_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AR_S13_HAS_SHRD_DDCTD_LNK
  `define AXI_AR_S13_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AR_S13_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AR_S13_NMV
  `define AXI_AR_S13_NMV `i_axi_AXI_AR_S13_NMV
`endif 

`ifdef i_axi_AXI_AR_S13_NMV_LOG2
  `define AXI_AR_S13_NMV_LOG2 `i_axi_AXI_AR_S13_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AR_S13_NMV_P1_LOG2
  `define AXI_AR_S13_NMV_P1_LOG2 `i_axi_AXI_AR_S13_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AW_S13_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AW_S13_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AW_S13_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AW_S13_HAS_SHRD_DDCTD_LNK
  `define AXI_AW_S13_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AW_S13_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AW_S13_NMV
  `define AXI_AW_S13_NMV `i_axi_AXI_AW_S13_NMV
`endif 

`ifdef i_axi_AXI_AW_S13_NMV_LOG2
  `define AXI_AW_S13_NMV_LOG2 `i_axi_AXI_AW_S13_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AW_S13_NMV_P1_LOG2
  `define AXI_AW_S13_NMV_P1_LOG2 `i_axi_AXI_AW_S13_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_W_S13_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_W_S13_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_W_S13_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_W_S13_HAS_SHRD_DDCTD_LNK
  `define AXI_W_S13_HAS_SHRD_DDCTD_LNK `i_axi_AXI_W_S13_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_W_S13_NMV
  `define AXI_W_S13_NMV `i_axi_AXI_W_S13_NMV
`endif 

`ifdef i_axi_AXI_W_S13_NMV_LOG2
  `define AXI_W_S13_NMV_LOG2 `i_axi_AXI_W_S13_NMV_LOG2
`endif 

`ifdef i_axi_AXI_W_S13_NMV_P1_LOG2
  `define AXI_W_S13_NMV_P1_LOG2 `i_axi_AXI_W_S13_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AR_S14_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AR_S14_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AR_S14_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AR_S14_HAS_SHRD_DDCTD_LNK
  `define AXI_AR_S14_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AR_S14_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AR_S14_NMV
  `define AXI_AR_S14_NMV `i_axi_AXI_AR_S14_NMV
`endif 

`ifdef i_axi_AXI_AR_S14_NMV_LOG2
  `define AXI_AR_S14_NMV_LOG2 `i_axi_AXI_AR_S14_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AR_S14_NMV_P1_LOG2
  `define AXI_AR_S14_NMV_P1_LOG2 `i_axi_AXI_AR_S14_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AW_S14_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AW_S14_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AW_S14_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AW_S14_HAS_SHRD_DDCTD_LNK
  `define AXI_AW_S14_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AW_S14_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AW_S14_NMV
  `define AXI_AW_S14_NMV `i_axi_AXI_AW_S14_NMV
`endif 

`ifdef i_axi_AXI_AW_S14_NMV_LOG2
  `define AXI_AW_S14_NMV_LOG2 `i_axi_AXI_AW_S14_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AW_S14_NMV_P1_LOG2
  `define AXI_AW_S14_NMV_P1_LOG2 `i_axi_AXI_AW_S14_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_W_S14_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_W_S14_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_W_S14_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_W_S14_HAS_SHRD_DDCTD_LNK
  `define AXI_W_S14_HAS_SHRD_DDCTD_LNK `i_axi_AXI_W_S14_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_W_S14_NMV
  `define AXI_W_S14_NMV `i_axi_AXI_W_S14_NMV
`endif 

`ifdef i_axi_AXI_W_S14_NMV_LOG2
  `define AXI_W_S14_NMV_LOG2 `i_axi_AXI_W_S14_NMV_LOG2
`endif 

`ifdef i_axi_AXI_W_S14_NMV_P1_LOG2
  `define AXI_W_S14_NMV_P1_LOG2 `i_axi_AXI_W_S14_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AR_S15_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AR_S15_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AR_S15_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AR_S15_HAS_SHRD_DDCTD_LNK
  `define AXI_AR_S15_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AR_S15_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AR_S15_NMV
  `define AXI_AR_S15_NMV `i_axi_AXI_AR_S15_NMV
`endif 

`ifdef i_axi_AXI_AR_S15_NMV_LOG2
  `define AXI_AR_S15_NMV_LOG2 `i_axi_AXI_AR_S15_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AR_S15_NMV_P1_LOG2
  `define AXI_AR_S15_NMV_P1_LOG2 `i_axi_AXI_AR_S15_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AW_S15_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AW_S15_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AW_S15_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AW_S15_HAS_SHRD_DDCTD_LNK
  `define AXI_AW_S15_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AW_S15_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AW_S15_NMV
  `define AXI_AW_S15_NMV `i_axi_AXI_AW_S15_NMV
`endif 

`ifdef i_axi_AXI_AW_S15_NMV_LOG2
  `define AXI_AW_S15_NMV_LOG2 `i_axi_AXI_AW_S15_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AW_S15_NMV_P1_LOG2
  `define AXI_AW_S15_NMV_P1_LOG2 `i_axi_AXI_AW_S15_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_W_S15_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_W_S15_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_W_S15_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_W_S15_HAS_SHRD_DDCTD_LNK
  `define AXI_W_S15_HAS_SHRD_DDCTD_LNK `i_axi_AXI_W_S15_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_W_S15_NMV
  `define AXI_W_S15_NMV `i_axi_AXI_W_S15_NMV
`endif 

`ifdef i_axi_AXI_W_S15_NMV_LOG2
  `define AXI_W_S15_NMV_LOG2 `i_axi_AXI_W_S15_NMV_LOG2
`endif 

`ifdef i_axi_AXI_W_S15_NMV_P1_LOG2
  `define AXI_W_S15_NMV_P1_LOG2 `i_axi_AXI_W_S15_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AR_S16_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AR_S16_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AR_S16_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AR_S16_HAS_SHRD_DDCTD_LNK
  `define AXI_AR_S16_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AR_S16_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AR_S16_NMV
  `define AXI_AR_S16_NMV `i_axi_AXI_AR_S16_NMV
`endif 

`ifdef i_axi_AXI_AR_S16_NMV_LOG2
  `define AXI_AR_S16_NMV_LOG2 `i_axi_AXI_AR_S16_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AR_S16_NMV_P1_LOG2
  `define AXI_AR_S16_NMV_P1_LOG2 `i_axi_AXI_AR_S16_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_AW_S16_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_AW_S16_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_AW_S16_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_AW_S16_HAS_SHRD_DDCTD_LNK
  `define AXI_AW_S16_HAS_SHRD_DDCTD_LNK `i_axi_AXI_AW_S16_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_AW_S16_NMV
  `define AXI_AW_S16_NMV `i_axi_AXI_AW_S16_NMV
`endif 

`ifdef i_axi_AXI_AW_S16_NMV_LOG2
  `define AXI_AW_S16_NMV_LOG2 `i_axi_AXI_AW_S16_NMV_LOG2
`endif 

`ifdef i_axi_AXI_AW_S16_NMV_P1_LOG2
  `define AXI_AW_S16_NMV_P1_LOG2 `i_axi_AXI_AW_S16_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_W_S16_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_W_S16_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_W_S16_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_W_S16_HAS_SHRD_DDCTD_LNK
  `define AXI_W_S16_HAS_SHRD_DDCTD_LNK `i_axi_AXI_W_S16_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_W_S16_NMV
  `define AXI_W_S16_NMV `i_axi_AXI_W_S16_NMV
`endif 

`ifdef i_axi_AXI_W_S16_NMV_LOG2
  `define AXI_W_S16_NMV_LOG2 `i_axi_AXI_W_S16_NMV_LOG2
`endif 

`ifdef i_axi_AXI_W_S16_NMV_P1_LOG2
  `define AXI_W_S16_NMV_P1_LOG2 `i_axi_AXI_W_S16_NMV_P1_LOG2
`endif 

`ifdef i_axi_AXI_R_M1_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_R_M1_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_R_M1_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_R_M1_HAS_SHRD_DDCTD_LNK
  `define AXI_R_M1_HAS_SHRD_DDCTD_LNK `i_axi_AXI_R_M1_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_R_M1_NSV
  `define AXI_R_M1_NSV `i_axi_AXI_R_M1_NSV
`endif 

`ifdef i_axi_AXI_R_M1_NSV_LOG2
  `define AXI_R_M1_NSV_LOG2 `i_axi_AXI_R_M1_NSV_LOG2
`endif 

`ifdef i_axi_AXI_R_M1_NSV_P1_LOG2
  `define AXI_R_M1_NSV_P1_LOG2 `i_axi_AXI_R_M1_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_B_M1_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_B_M1_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_B_M1_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_B_M1_HAS_SHRD_DDCTD_LNK
  `define AXI_B_M1_HAS_SHRD_DDCTD_LNK `i_axi_AXI_B_M1_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_B_M1_NSV
  `define AXI_B_M1_NSV `i_axi_AXI_B_M1_NSV
`endif 

`ifdef i_axi_AXI_B_M1_NSV_LOG2
  `define AXI_B_M1_NSV_LOG2 `i_axi_AXI_B_M1_NSV_LOG2
`endif 

`ifdef i_axi_AXI_B_M1_NSV_P1_LOG2
  `define AXI_B_M1_NSV_P1_LOG2 `i_axi_AXI_B_M1_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_R_M2_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_R_M2_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_R_M2_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_R_M2_HAS_SHRD_DDCTD_LNK
  `define AXI_R_M2_HAS_SHRD_DDCTD_LNK `i_axi_AXI_R_M2_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_R_M2_NSV
  `define AXI_R_M2_NSV `i_axi_AXI_R_M2_NSV
`endif 

`ifdef i_axi_AXI_R_M2_NSV_LOG2
  `define AXI_R_M2_NSV_LOG2 `i_axi_AXI_R_M2_NSV_LOG2
`endif 

`ifdef i_axi_AXI_R_M2_NSV_P1_LOG2
  `define AXI_R_M2_NSV_P1_LOG2 `i_axi_AXI_R_M2_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_B_M2_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_B_M2_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_B_M2_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_B_M2_HAS_SHRD_DDCTD_LNK
  `define AXI_B_M2_HAS_SHRD_DDCTD_LNK `i_axi_AXI_B_M2_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_B_M2_NSV
  `define AXI_B_M2_NSV `i_axi_AXI_B_M2_NSV
`endif 

`ifdef i_axi_AXI_B_M2_NSV_LOG2
  `define AXI_B_M2_NSV_LOG2 `i_axi_AXI_B_M2_NSV_LOG2
`endif 

`ifdef i_axi_AXI_B_M2_NSV_P1_LOG2
  `define AXI_B_M2_NSV_P1_LOG2 `i_axi_AXI_B_M2_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_R_M3_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_R_M3_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_R_M3_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_R_M3_HAS_SHRD_DDCTD_LNK
  `define AXI_R_M3_HAS_SHRD_DDCTD_LNK `i_axi_AXI_R_M3_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_R_M3_NSV
  `define AXI_R_M3_NSV `i_axi_AXI_R_M3_NSV
`endif 

`ifdef i_axi_AXI_R_M3_NSV_LOG2
  `define AXI_R_M3_NSV_LOG2 `i_axi_AXI_R_M3_NSV_LOG2
`endif 

`ifdef i_axi_AXI_R_M3_NSV_P1_LOG2
  `define AXI_R_M3_NSV_P1_LOG2 `i_axi_AXI_R_M3_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_B_M3_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_B_M3_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_B_M3_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_B_M3_HAS_SHRD_DDCTD_LNK
  `define AXI_B_M3_HAS_SHRD_DDCTD_LNK `i_axi_AXI_B_M3_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_B_M3_NSV
  `define AXI_B_M3_NSV `i_axi_AXI_B_M3_NSV
`endif 

`ifdef i_axi_AXI_B_M3_NSV_LOG2
  `define AXI_B_M3_NSV_LOG2 `i_axi_AXI_B_M3_NSV_LOG2
`endif 

`ifdef i_axi_AXI_B_M3_NSV_P1_LOG2
  `define AXI_B_M3_NSV_P1_LOG2 `i_axi_AXI_B_M3_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_R_M4_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_R_M4_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_R_M4_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_R_M4_HAS_SHRD_DDCTD_LNK
  `define AXI_R_M4_HAS_SHRD_DDCTD_LNK `i_axi_AXI_R_M4_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_R_M4_NSV
  `define AXI_R_M4_NSV `i_axi_AXI_R_M4_NSV
`endif 

`ifdef i_axi_AXI_R_M4_NSV_LOG2
  `define AXI_R_M4_NSV_LOG2 `i_axi_AXI_R_M4_NSV_LOG2
`endif 

`ifdef i_axi_AXI_R_M4_NSV_P1_LOG2
  `define AXI_R_M4_NSV_P1_LOG2 `i_axi_AXI_R_M4_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_B_M4_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_B_M4_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_B_M4_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_B_M4_HAS_SHRD_DDCTD_LNK
  `define AXI_B_M4_HAS_SHRD_DDCTD_LNK `i_axi_AXI_B_M4_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_B_M4_NSV
  `define AXI_B_M4_NSV `i_axi_AXI_B_M4_NSV
`endif 

`ifdef i_axi_AXI_B_M4_NSV_LOG2
  `define AXI_B_M4_NSV_LOG2 `i_axi_AXI_B_M4_NSV_LOG2
`endif 

`ifdef i_axi_AXI_B_M4_NSV_P1_LOG2
  `define AXI_B_M4_NSV_P1_LOG2 `i_axi_AXI_B_M4_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_R_M5_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_R_M5_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_R_M5_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_R_M5_HAS_SHRD_DDCTD_LNK
  `define AXI_R_M5_HAS_SHRD_DDCTD_LNK `i_axi_AXI_R_M5_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_R_M5_NSV
  `define AXI_R_M5_NSV `i_axi_AXI_R_M5_NSV
`endif 

`ifdef i_axi_AXI_R_M5_NSV_LOG2
  `define AXI_R_M5_NSV_LOG2 `i_axi_AXI_R_M5_NSV_LOG2
`endif 

`ifdef i_axi_AXI_R_M5_NSV_P1_LOG2
  `define AXI_R_M5_NSV_P1_LOG2 `i_axi_AXI_R_M5_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_B_M5_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_B_M5_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_B_M5_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_B_M5_HAS_SHRD_DDCTD_LNK
  `define AXI_B_M5_HAS_SHRD_DDCTD_LNK `i_axi_AXI_B_M5_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_B_M5_NSV
  `define AXI_B_M5_NSV `i_axi_AXI_B_M5_NSV
`endif 

`ifdef i_axi_AXI_B_M5_NSV_LOG2
  `define AXI_B_M5_NSV_LOG2 `i_axi_AXI_B_M5_NSV_LOG2
`endif 

`ifdef i_axi_AXI_B_M5_NSV_P1_LOG2
  `define AXI_B_M5_NSV_P1_LOG2 `i_axi_AXI_B_M5_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_R_M6_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_R_M6_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_R_M6_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_R_M6_HAS_SHRD_DDCTD_LNK
  `define AXI_R_M6_HAS_SHRD_DDCTD_LNK `i_axi_AXI_R_M6_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_R_M6_NSV
  `define AXI_R_M6_NSV `i_axi_AXI_R_M6_NSV
`endif 

`ifdef i_axi_AXI_R_M6_NSV_LOG2
  `define AXI_R_M6_NSV_LOG2 `i_axi_AXI_R_M6_NSV_LOG2
`endif 

`ifdef i_axi_AXI_R_M6_NSV_P1_LOG2
  `define AXI_R_M6_NSV_P1_LOG2 `i_axi_AXI_R_M6_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_B_M6_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_B_M6_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_B_M6_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_B_M6_HAS_SHRD_DDCTD_LNK
  `define AXI_B_M6_HAS_SHRD_DDCTD_LNK `i_axi_AXI_B_M6_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_B_M6_NSV
  `define AXI_B_M6_NSV `i_axi_AXI_B_M6_NSV
`endif 

`ifdef i_axi_AXI_B_M6_NSV_LOG2
  `define AXI_B_M6_NSV_LOG2 `i_axi_AXI_B_M6_NSV_LOG2
`endif 

`ifdef i_axi_AXI_B_M6_NSV_P1_LOG2
  `define AXI_B_M6_NSV_P1_LOG2 `i_axi_AXI_B_M6_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_R_M7_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_R_M7_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_R_M7_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_R_M7_HAS_SHRD_DDCTD_LNK
  `define AXI_R_M7_HAS_SHRD_DDCTD_LNK `i_axi_AXI_R_M7_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_R_M7_NSV
  `define AXI_R_M7_NSV `i_axi_AXI_R_M7_NSV
`endif 

`ifdef i_axi_AXI_R_M7_NSV_LOG2
  `define AXI_R_M7_NSV_LOG2 `i_axi_AXI_R_M7_NSV_LOG2
`endif 

`ifdef i_axi_AXI_R_M7_NSV_P1_LOG2
  `define AXI_R_M7_NSV_P1_LOG2 `i_axi_AXI_R_M7_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_B_M7_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_B_M7_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_B_M7_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_B_M7_HAS_SHRD_DDCTD_LNK
  `define AXI_B_M7_HAS_SHRD_DDCTD_LNK `i_axi_AXI_B_M7_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_B_M7_NSV
  `define AXI_B_M7_NSV `i_axi_AXI_B_M7_NSV
`endif 

`ifdef i_axi_AXI_B_M7_NSV_LOG2
  `define AXI_B_M7_NSV_LOG2 `i_axi_AXI_B_M7_NSV_LOG2
`endif 

`ifdef i_axi_AXI_B_M7_NSV_P1_LOG2
  `define AXI_B_M7_NSV_P1_LOG2 `i_axi_AXI_B_M7_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_R_M8_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_R_M8_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_R_M8_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_R_M8_HAS_SHRD_DDCTD_LNK
  `define AXI_R_M8_HAS_SHRD_DDCTD_LNK `i_axi_AXI_R_M8_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_R_M8_NSV
  `define AXI_R_M8_NSV `i_axi_AXI_R_M8_NSV
`endif 

`ifdef i_axi_AXI_R_M8_NSV_LOG2
  `define AXI_R_M8_NSV_LOG2 `i_axi_AXI_R_M8_NSV_LOG2
`endif 

`ifdef i_axi_AXI_R_M8_NSV_P1_LOG2
  `define AXI_R_M8_NSV_P1_LOG2 `i_axi_AXI_R_M8_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_B_M8_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_B_M8_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_B_M8_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_B_M8_HAS_SHRD_DDCTD_LNK
  `define AXI_B_M8_HAS_SHRD_DDCTD_LNK `i_axi_AXI_B_M8_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_B_M8_NSV
  `define AXI_B_M8_NSV `i_axi_AXI_B_M8_NSV
`endif 

`ifdef i_axi_AXI_B_M8_NSV_LOG2
  `define AXI_B_M8_NSV_LOG2 `i_axi_AXI_B_M8_NSV_LOG2
`endif 

`ifdef i_axi_AXI_B_M8_NSV_P1_LOG2
  `define AXI_B_M8_NSV_P1_LOG2 `i_axi_AXI_B_M8_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_R_M9_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_R_M9_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_R_M9_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_R_M9_HAS_SHRD_DDCTD_LNK
  `define AXI_R_M9_HAS_SHRD_DDCTD_LNK `i_axi_AXI_R_M9_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_R_M9_NSV
  `define AXI_R_M9_NSV `i_axi_AXI_R_M9_NSV
`endif 

`ifdef i_axi_AXI_R_M9_NSV_LOG2
  `define AXI_R_M9_NSV_LOG2 `i_axi_AXI_R_M9_NSV_LOG2
`endif 

`ifdef i_axi_AXI_R_M9_NSV_P1_LOG2
  `define AXI_R_M9_NSV_P1_LOG2 `i_axi_AXI_R_M9_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_B_M9_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_B_M9_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_B_M9_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_B_M9_HAS_SHRD_DDCTD_LNK
  `define AXI_B_M9_HAS_SHRD_DDCTD_LNK `i_axi_AXI_B_M9_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_B_M9_NSV
  `define AXI_B_M9_NSV `i_axi_AXI_B_M9_NSV
`endif 

`ifdef i_axi_AXI_B_M9_NSV_LOG2
  `define AXI_B_M9_NSV_LOG2 `i_axi_AXI_B_M9_NSV_LOG2
`endif 

`ifdef i_axi_AXI_B_M9_NSV_P1_LOG2
  `define AXI_B_M9_NSV_P1_LOG2 `i_axi_AXI_B_M9_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_R_M10_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_R_M10_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_R_M10_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_R_M10_HAS_SHRD_DDCTD_LNK
  `define AXI_R_M10_HAS_SHRD_DDCTD_LNK `i_axi_AXI_R_M10_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_R_M10_NSV
  `define AXI_R_M10_NSV `i_axi_AXI_R_M10_NSV
`endif 

`ifdef i_axi_AXI_R_M10_NSV_LOG2
  `define AXI_R_M10_NSV_LOG2 `i_axi_AXI_R_M10_NSV_LOG2
`endif 

`ifdef i_axi_AXI_R_M10_NSV_P1_LOG2
  `define AXI_R_M10_NSV_P1_LOG2 `i_axi_AXI_R_M10_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_B_M10_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_B_M10_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_B_M10_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_B_M10_HAS_SHRD_DDCTD_LNK
  `define AXI_B_M10_HAS_SHRD_DDCTD_LNK `i_axi_AXI_B_M10_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_B_M10_NSV
  `define AXI_B_M10_NSV `i_axi_AXI_B_M10_NSV
`endif 

`ifdef i_axi_AXI_B_M10_NSV_LOG2
  `define AXI_B_M10_NSV_LOG2 `i_axi_AXI_B_M10_NSV_LOG2
`endif 

`ifdef i_axi_AXI_B_M10_NSV_P1_LOG2
  `define AXI_B_M10_NSV_P1_LOG2 `i_axi_AXI_B_M10_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_R_M11_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_R_M11_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_R_M11_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_R_M11_HAS_SHRD_DDCTD_LNK
  `define AXI_R_M11_HAS_SHRD_DDCTD_LNK `i_axi_AXI_R_M11_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_R_M11_NSV
  `define AXI_R_M11_NSV `i_axi_AXI_R_M11_NSV
`endif 

`ifdef i_axi_AXI_R_M11_NSV_LOG2
  `define AXI_R_M11_NSV_LOG2 `i_axi_AXI_R_M11_NSV_LOG2
`endif 

`ifdef i_axi_AXI_R_M11_NSV_P1_LOG2
  `define AXI_R_M11_NSV_P1_LOG2 `i_axi_AXI_R_M11_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_B_M11_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_B_M11_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_B_M11_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_B_M11_HAS_SHRD_DDCTD_LNK
  `define AXI_B_M11_HAS_SHRD_DDCTD_LNK `i_axi_AXI_B_M11_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_B_M11_NSV
  `define AXI_B_M11_NSV `i_axi_AXI_B_M11_NSV
`endif 

`ifdef i_axi_AXI_B_M11_NSV_LOG2
  `define AXI_B_M11_NSV_LOG2 `i_axi_AXI_B_M11_NSV_LOG2
`endif 

`ifdef i_axi_AXI_B_M11_NSV_P1_LOG2
  `define AXI_B_M11_NSV_P1_LOG2 `i_axi_AXI_B_M11_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_R_M12_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_R_M12_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_R_M12_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_R_M12_HAS_SHRD_DDCTD_LNK
  `define AXI_R_M12_HAS_SHRD_DDCTD_LNK `i_axi_AXI_R_M12_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_R_M12_NSV
  `define AXI_R_M12_NSV `i_axi_AXI_R_M12_NSV
`endif 

`ifdef i_axi_AXI_R_M12_NSV_LOG2
  `define AXI_R_M12_NSV_LOG2 `i_axi_AXI_R_M12_NSV_LOG2
`endif 

`ifdef i_axi_AXI_R_M12_NSV_P1_LOG2
  `define AXI_R_M12_NSV_P1_LOG2 `i_axi_AXI_R_M12_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_B_M12_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_B_M12_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_B_M12_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_B_M12_HAS_SHRD_DDCTD_LNK
  `define AXI_B_M12_HAS_SHRD_DDCTD_LNK `i_axi_AXI_B_M12_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_B_M12_NSV
  `define AXI_B_M12_NSV `i_axi_AXI_B_M12_NSV
`endif 

`ifdef i_axi_AXI_B_M12_NSV_LOG2
  `define AXI_B_M12_NSV_LOG2 `i_axi_AXI_B_M12_NSV_LOG2
`endif 

`ifdef i_axi_AXI_B_M12_NSV_P1_LOG2
  `define AXI_B_M12_NSV_P1_LOG2 `i_axi_AXI_B_M12_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_R_M13_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_R_M13_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_R_M13_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_R_M13_HAS_SHRD_DDCTD_LNK
  `define AXI_R_M13_HAS_SHRD_DDCTD_LNK `i_axi_AXI_R_M13_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_R_M13_NSV
  `define AXI_R_M13_NSV `i_axi_AXI_R_M13_NSV
`endif 

`ifdef i_axi_AXI_R_M13_NSV_LOG2
  `define AXI_R_M13_NSV_LOG2 `i_axi_AXI_R_M13_NSV_LOG2
`endif 

`ifdef i_axi_AXI_R_M13_NSV_P1_LOG2
  `define AXI_R_M13_NSV_P1_LOG2 `i_axi_AXI_R_M13_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_B_M13_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_B_M13_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_B_M13_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_B_M13_HAS_SHRD_DDCTD_LNK
  `define AXI_B_M13_HAS_SHRD_DDCTD_LNK `i_axi_AXI_B_M13_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_B_M13_NSV
  `define AXI_B_M13_NSV `i_axi_AXI_B_M13_NSV
`endif 

`ifdef i_axi_AXI_B_M13_NSV_LOG2
  `define AXI_B_M13_NSV_LOG2 `i_axi_AXI_B_M13_NSV_LOG2
`endif 

`ifdef i_axi_AXI_B_M13_NSV_P1_LOG2
  `define AXI_B_M13_NSV_P1_LOG2 `i_axi_AXI_B_M13_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_R_M14_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_R_M14_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_R_M14_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_R_M14_HAS_SHRD_DDCTD_LNK
  `define AXI_R_M14_HAS_SHRD_DDCTD_LNK `i_axi_AXI_R_M14_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_R_M14_NSV
  `define AXI_R_M14_NSV `i_axi_AXI_R_M14_NSV
`endif 

`ifdef i_axi_AXI_R_M14_NSV_LOG2
  `define AXI_R_M14_NSV_LOG2 `i_axi_AXI_R_M14_NSV_LOG2
`endif 

`ifdef i_axi_AXI_R_M14_NSV_P1_LOG2
  `define AXI_R_M14_NSV_P1_LOG2 `i_axi_AXI_R_M14_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_B_M14_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_B_M14_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_B_M14_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_B_M14_HAS_SHRD_DDCTD_LNK
  `define AXI_B_M14_HAS_SHRD_DDCTD_LNK `i_axi_AXI_B_M14_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_B_M14_NSV
  `define AXI_B_M14_NSV `i_axi_AXI_B_M14_NSV
`endif 

`ifdef i_axi_AXI_B_M14_NSV_LOG2
  `define AXI_B_M14_NSV_LOG2 `i_axi_AXI_B_M14_NSV_LOG2
`endif 

`ifdef i_axi_AXI_B_M14_NSV_P1_LOG2
  `define AXI_B_M14_NSV_P1_LOG2 `i_axi_AXI_B_M14_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_R_M15_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_R_M15_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_R_M15_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_R_M15_HAS_SHRD_DDCTD_LNK
  `define AXI_R_M15_HAS_SHRD_DDCTD_LNK `i_axi_AXI_R_M15_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_R_M15_NSV
  `define AXI_R_M15_NSV `i_axi_AXI_R_M15_NSV
`endif 

`ifdef i_axi_AXI_R_M15_NSV_LOG2
  `define AXI_R_M15_NSV_LOG2 `i_axi_AXI_R_M15_NSV_LOG2
`endif 

`ifdef i_axi_AXI_R_M15_NSV_P1_LOG2
  `define AXI_R_M15_NSV_P1_LOG2 `i_axi_AXI_R_M15_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_B_M15_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_B_M15_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_B_M15_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_B_M15_HAS_SHRD_DDCTD_LNK
  `define AXI_B_M15_HAS_SHRD_DDCTD_LNK `i_axi_AXI_B_M15_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_B_M15_NSV
  `define AXI_B_M15_NSV `i_axi_AXI_B_M15_NSV
`endif 

`ifdef i_axi_AXI_B_M15_NSV_LOG2
  `define AXI_B_M15_NSV_LOG2 `i_axi_AXI_B_M15_NSV_LOG2
`endif 

`ifdef i_axi_AXI_B_M15_NSV_P1_LOG2
  `define AXI_B_M15_NSV_P1_LOG2 `i_axi_AXI_B_M15_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_R_M16_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_R_M16_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_R_M16_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_R_M16_HAS_SHRD_DDCTD_LNK
  `define AXI_R_M16_HAS_SHRD_DDCTD_LNK `i_axi_AXI_R_M16_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_R_M16_NSV
  `define AXI_R_M16_NSV `i_axi_AXI_R_M16_NSV
`endif 

`ifdef i_axi_AXI_R_M16_NSV_LOG2
  `define AXI_R_M16_NSV_LOG2 `i_axi_AXI_R_M16_NSV_LOG2
`endif 

`ifdef i_axi_AXI_R_M16_NSV_P1_LOG2
  `define AXI_R_M16_NSV_P1_LOG2 `i_axi_AXI_R_M16_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_B_M16_HAS_SHRD_DDCTD_LNK_VAL
  `define AXI_B_M16_HAS_SHRD_DDCTD_LNK_VAL `i_axi_AXI_B_M16_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef i_axi_AXI_B_M16_HAS_SHRD_DDCTD_LNK
  `define AXI_B_M16_HAS_SHRD_DDCTD_LNK `i_axi_AXI_B_M16_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef i_axi_AXI_B_M16_NSV
  `define AXI_B_M16_NSV `i_axi_AXI_B_M16_NSV
`endif 

`ifdef i_axi_AXI_B_M16_NSV_LOG2
  `define AXI_B_M16_NSV_LOG2 `i_axi_AXI_B_M16_NSV_LOG2
`endif 

`ifdef i_axi_AXI_B_M16_NSV_P1_LOG2
  `define AXI_B_M16_NSV_P1_LOG2 `i_axi_AXI_B_M16_NSV_P1_LOG2
`endif 

`ifdef i_axi_AXI_M1_ON_AR_SHARED_VAL
  `define AXI_M1_ON_AR_SHARED_VAL `i_axi_AXI_M1_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M2_ON_AR_SHARED_VAL
  `define AXI_M2_ON_AR_SHARED_VAL `i_axi_AXI_M2_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M3_ON_AR_SHARED_VAL
  `define AXI_M3_ON_AR_SHARED_VAL `i_axi_AXI_M3_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M4_ON_AR_SHARED_VAL
  `define AXI_M4_ON_AR_SHARED_VAL `i_axi_AXI_M4_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M5_ON_AR_SHARED_VAL
  `define AXI_M5_ON_AR_SHARED_VAL `i_axi_AXI_M5_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M6_ON_AR_SHARED_VAL
  `define AXI_M6_ON_AR_SHARED_VAL `i_axi_AXI_M6_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M7_ON_AR_SHARED_VAL
  `define AXI_M7_ON_AR_SHARED_VAL `i_axi_AXI_M7_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M8_ON_AR_SHARED_VAL
  `define AXI_M8_ON_AR_SHARED_VAL `i_axi_AXI_M8_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M9_ON_AR_SHARED_VAL
  `define AXI_M9_ON_AR_SHARED_VAL `i_axi_AXI_M9_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M10_ON_AR_SHARED_VAL
  `define AXI_M10_ON_AR_SHARED_VAL `i_axi_AXI_M10_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M11_ON_AR_SHARED_VAL
  `define AXI_M11_ON_AR_SHARED_VAL `i_axi_AXI_M11_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M12_ON_AR_SHARED_VAL
  `define AXI_M12_ON_AR_SHARED_VAL `i_axi_AXI_M12_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M13_ON_AR_SHARED_VAL
  `define AXI_M13_ON_AR_SHARED_VAL `i_axi_AXI_M13_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M14_ON_AR_SHARED_VAL
  `define AXI_M14_ON_AR_SHARED_VAL `i_axi_AXI_M14_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M15_ON_AR_SHARED_VAL
  `define AXI_M15_ON_AR_SHARED_VAL `i_axi_AXI_M15_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M16_ON_AR_SHARED_VAL
  `define AXI_M16_ON_AR_SHARED_VAL `i_axi_AXI_M16_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S0_ON_AR_SHARED_VAL
  `define AXI_S0_ON_AR_SHARED_VAL `i_axi_AXI_S0_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S0_ON_AR_SHARED_ONLY
  `define AXI_S0_ON_AR_SHARED_ONLY `i_axi_AXI_S0_ON_AR_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S0_ON_AR_SHARED_ONLY_VAL
  `define AXI_S0_ON_AR_SHARED_ONLY_VAL `i_axi_AXI_S0_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S1_ON_AR_SHARED_VAL
  `define AXI_S1_ON_AR_SHARED_VAL `i_axi_AXI_S1_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S1_ON_AR_SHARED_ONLY
  `define AXI_S1_ON_AR_SHARED_ONLY `i_axi_AXI_S1_ON_AR_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S1_ON_AR_SHARED_ONLY_VAL
  `define AXI_S1_ON_AR_SHARED_ONLY_VAL `i_axi_AXI_S1_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S2_ON_AR_SHARED_VAL
  `define AXI_S2_ON_AR_SHARED_VAL `i_axi_AXI_S2_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S2_ON_AR_SHARED_ONLY
  `define AXI_S2_ON_AR_SHARED_ONLY `i_axi_AXI_S2_ON_AR_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S2_ON_AR_SHARED_ONLY_VAL
  `define AXI_S2_ON_AR_SHARED_ONLY_VAL `i_axi_AXI_S2_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S3_ON_AR_SHARED_VAL
  `define AXI_S3_ON_AR_SHARED_VAL `i_axi_AXI_S3_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S3_ON_AR_SHARED_ONLY
  `define AXI_S3_ON_AR_SHARED_ONLY `i_axi_AXI_S3_ON_AR_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S3_ON_AR_SHARED_ONLY_VAL
  `define AXI_S3_ON_AR_SHARED_ONLY_VAL `i_axi_AXI_S3_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S4_ON_AR_SHARED_VAL
  `define AXI_S4_ON_AR_SHARED_VAL `i_axi_AXI_S4_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S4_ON_AR_SHARED_ONLY
  `define AXI_S4_ON_AR_SHARED_ONLY `i_axi_AXI_S4_ON_AR_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S4_ON_AR_SHARED_ONLY_VAL
  `define AXI_S4_ON_AR_SHARED_ONLY_VAL `i_axi_AXI_S4_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S5_ON_AR_SHARED_VAL
  `define AXI_S5_ON_AR_SHARED_VAL `i_axi_AXI_S5_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S5_ON_AR_SHARED_ONLY
  `define AXI_S5_ON_AR_SHARED_ONLY `i_axi_AXI_S5_ON_AR_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S5_ON_AR_SHARED_ONLY_VAL
  `define AXI_S5_ON_AR_SHARED_ONLY_VAL `i_axi_AXI_S5_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S6_ON_AR_SHARED_VAL
  `define AXI_S6_ON_AR_SHARED_VAL `i_axi_AXI_S6_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S6_ON_AR_SHARED_ONLY
  `define AXI_S6_ON_AR_SHARED_ONLY `i_axi_AXI_S6_ON_AR_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S6_ON_AR_SHARED_ONLY_VAL
  `define AXI_S6_ON_AR_SHARED_ONLY_VAL `i_axi_AXI_S6_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S7_ON_AR_SHARED_VAL
  `define AXI_S7_ON_AR_SHARED_VAL `i_axi_AXI_S7_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S7_ON_AR_SHARED_ONLY
  `define AXI_S7_ON_AR_SHARED_ONLY `i_axi_AXI_S7_ON_AR_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S7_ON_AR_SHARED_ONLY_VAL
  `define AXI_S7_ON_AR_SHARED_ONLY_VAL `i_axi_AXI_S7_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S8_ON_AR_SHARED_VAL
  `define AXI_S8_ON_AR_SHARED_VAL `i_axi_AXI_S8_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S8_ON_AR_SHARED_ONLY
  `define AXI_S8_ON_AR_SHARED_ONLY `i_axi_AXI_S8_ON_AR_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S8_ON_AR_SHARED_ONLY_VAL
  `define AXI_S8_ON_AR_SHARED_ONLY_VAL `i_axi_AXI_S8_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S9_ON_AR_SHARED_VAL
  `define AXI_S9_ON_AR_SHARED_VAL `i_axi_AXI_S9_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S9_ON_AR_SHARED_ONLY
  `define AXI_S9_ON_AR_SHARED_ONLY `i_axi_AXI_S9_ON_AR_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S9_ON_AR_SHARED_ONLY_VAL
  `define AXI_S9_ON_AR_SHARED_ONLY_VAL `i_axi_AXI_S9_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S10_ON_AR_SHARED_VAL
  `define AXI_S10_ON_AR_SHARED_VAL `i_axi_AXI_S10_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S10_ON_AR_SHARED_ONLY
  `define AXI_S10_ON_AR_SHARED_ONLY `i_axi_AXI_S10_ON_AR_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S10_ON_AR_SHARED_ONLY_VAL
  `define AXI_S10_ON_AR_SHARED_ONLY_VAL `i_axi_AXI_S10_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S11_ON_AR_SHARED_VAL
  `define AXI_S11_ON_AR_SHARED_VAL `i_axi_AXI_S11_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S11_ON_AR_SHARED_ONLY
  `define AXI_S11_ON_AR_SHARED_ONLY `i_axi_AXI_S11_ON_AR_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S11_ON_AR_SHARED_ONLY_VAL
  `define AXI_S11_ON_AR_SHARED_ONLY_VAL `i_axi_AXI_S11_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S12_ON_AR_SHARED_VAL
  `define AXI_S12_ON_AR_SHARED_VAL `i_axi_AXI_S12_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S12_ON_AR_SHARED_ONLY
  `define AXI_S12_ON_AR_SHARED_ONLY `i_axi_AXI_S12_ON_AR_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S12_ON_AR_SHARED_ONLY_VAL
  `define AXI_S12_ON_AR_SHARED_ONLY_VAL `i_axi_AXI_S12_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S13_ON_AR_SHARED_VAL
  `define AXI_S13_ON_AR_SHARED_VAL `i_axi_AXI_S13_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S13_ON_AR_SHARED_ONLY
  `define AXI_S13_ON_AR_SHARED_ONLY `i_axi_AXI_S13_ON_AR_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S13_ON_AR_SHARED_ONLY_VAL
  `define AXI_S13_ON_AR_SHARED_ONLY_VAL `i_axi_AXI_S13_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S14_ON_AR_SHARED_VAL
  `define AXI_S14_ON_AR_SHARED_VAL `i_axi_AXI_S14_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S14_ON_AR_SHARED_ONLY
  `define AXI_S14_ON_AR_SHARED_ONLY `i_axi_AXI_S14_ON_AR_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S14_ON_AR_SHARED_ONLY_VAL
  `define AXI_S14_ON_AR_SHARED_ONLY_VAL `i_axi_AXI_S14_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S15_ON_AR_SHARED_VAL
  `define AXI_S15_ON_AR_SHARED_VAL `i_axi_AXI_S15_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S15_ON_AR_SHARED_ONLY
  `define AXI_S15_ON_AR_SHARED_ONLY `i_axi_AXI_S15_ON_AR_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S15_ON_AR_SHARED_ONLY_VAL
  `define AXI_S15_ON_AR_SHARED_ONLY_VAL `i_axi_AXI_S15_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S16_ON_AR_SHARED_VAL
  `define AXI_S16_ON_AR_SHARED_VAL `i_axi_AXI_S16_ON_AR_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S16_ON_AR_SHARED_ONLY
  `define AXI_S16_ON_AR_SHARED_ONLY `i_axi_AXI_S16_ON_AR_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S16_ON_AR_SHARED_ONLY_VAL
  `define AXI_S16_ON_AR_SHARED_ONLY_VAL `i_axi_AXI_S16_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M1_ON_AW_SHARED_VAL
  `define AXI_M1_ON_AW_SHARED_VAL `i_axi_AXI_M1_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M2_ON_AW_SHARED_VAL
  `define AXI_M2_ON_AW_SHARED_VAL `i_axi_AXI_M2_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M3_ON_AW_SHARED_VAL
  `define AXI_M3_ON_AW_SHARED_VAL `i_axi_AXI_M3_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M4_ON_AW_SHARED_VAL
  `define AXI_M4_ON_AW_SHARED_VAL `i_axi_AXI_M4_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M5_ON_AW_SHARED_VAL
  `define AXI_M5_ON_AW_SHARED_VAL `i_axi_AXI_M5_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M6_ON_AW_SHARED_VAL
  `define AXI_M6_ON_AW_SHARED_VAL `i_axi_AXI_M6_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M7_ON_AW_SHARED_VAL
  `define AXI_M7_ON_AW_SHARED_VAL `i_axi_AXI_M7_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M8_ON_AW_SHARED_VAL
  `define AXI_M8_ON_AW_SHARED_VAL `i_axi_AXI_M8_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M9_ON_AW_SHARED_VAL
  `define AXI_M9_ON_AW_SHARED_VAL `i_axi_AXI_M9_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M10_ON_AW_SHARED_VAL
  `define AXI_M10_ON_AW_SHARED_VAL `i_axi_AXI_M10_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M11_ON_AW_SHARED_VAL
  `define AXI_M11_ON_AW_SHARED_VAL `i_axi_AXI_M11_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M12_ON_AW_SHARED_VAL
  `define AXI_M12_ON_AW_SHARED_VAL `i_axi_AXI_M12_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M13_ON_AW_SHARED_VAL
  `define AXI_M13_ON_AW_SHARED_VAL `i_axi_AXI_M13_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M14_ON_AW_SHARED_VAL
  `define AXI_M14_ON_AW_SHARED_VAL `i_axi_AXI_M14_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M15_ON_AW_SHARED_VAL
  `define AXI_M15_ON_AW_SHARED_VAL `i_axi_AXI_M15_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M16_ON_AW_SHARED_VAL
  `define AXI_M16_ON_AW_SHARED_VAL `i_axi_AXI_M16_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S0_ON_AW_SHARED_VAL
  `define AXI_S0_ON_AW_SHARED_VAL `i_axi_AXI_S0_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S0_ON_AW_SHARED_ONLY
  `define AXI_S0_ON_AW_SHARED_ONLY `i_axi_AXI_S0_ON_AW_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S0_ON_AW_SHARED_ONLY_VAL
  `define AXI_S0_ON_AW_SHARED_ONLY_VAL `i_axi_AXI_S0_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S1_ON_AW_SHARED_VAL
  `define AXI_S1_ON_AW_SHARED_VAL `i_axi_AXI_S1_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S1_ON_AW_SHARED_ONLY
  `define AXI_S1_ON_AW_SHARED_ONLY `i_axi_AXI_S1_ON_AW_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S1_ON_AW_SHARED_ONLY_VAL
  `define AXI_S1_ON_AW_SHARED_ONLY_VAL `i_axi_AXI_S1_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S2_ON_AW_SHARED_VAL
  `define AXI_S2_ON_AW_SHARED_VAL `i_axi_AXI_S2_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S2_ON_AW_SHARED_ONLY
  `define AXI_S2_ON_AW_SHARED_ONLY `i_axi_AXI_S2_ON_AW_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S2_ON_AW_SHARED_ONLY_VAL
  `define AXI_S2_ON_AW_SHARED_ONLY_VAL `i_axi_AXI_S2_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S3_ON_AW_SHARED_VAL
  `define AXI_S3_ON_AW_SHARED_VAL `i_axi_AXI_S3_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S3_ON_AW_SHARED_ONLY
  `define AXI_S3_ON_AW_SHARED_ONLY `i_axi_AXI_S3_ON_AW_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S3_ON_AW_SHARED_ONLY_VAL
  `define AXI_S3_ON_AW_SHARED_ONLY_VAL `i_axi_AXI_S3_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S4_ON_AW_SHARED_VAL
  `define AXI_S4_ON_AW_SHARED_VAL `i_axi_AXI_S4_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S4_ON_AW_SHARED_ONLY
  `define AXI_S4_ON_AW_SHARED_ONLY `i_axi_AXI_S4_ON_AW_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S4_ON_AW_SHARED_ONLY_VAL
  `define AXI_S4_ON_AW_SHARED_ONLY_VAL `i_axi_AXI_S4_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S5_ON_AW_SHARED_VAL
  `define AXI_S5_ON_AW_SHARED_VAL `i_axi_AXI_S5_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S5_ON_AW_SHARED_ONLY
  `define AXI_S5_ON_AW_SHARED_ONLY `i_axi_AXI_S5_ON_AW_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S5_ON_AW_SHARED_ONLY_VAL
  `define AXI_S5_ON_AW_SHARED_ONLY_VAL `i_axi_AXI_S5_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S6_ON_AW_SHARED_VAL
  `define AXI_S6_ON_AW_SHARED_VAL `i_axi_AXI_S6_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S6_ON_AW_SHARED_ONLY
  `define AXI_S6_ON_AW_SHARED_ONLY `i_axi_AXI_S6_ON_AW_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S6_ON_AW_SHARED_ONLY_VAL
  `define AXI_S6_ON_AW_SHARED_ONLY_VAL `i_axi_AXI_S6_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S7_ON_AW_SHARED_VAL
  `define AXI_S7_ON_AW_SHARED_VAL `i_axi_AXI_S7_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S7_ON_AW_SHARED_ONLY
  `define AXI_S7_ON_AW_SHARED_ONLY `i_axi_AXI_S7_ON_AW_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S7_ON_AW_SHARED_ONLY_VAL
  `define AXI_S7_ON_AW_SHARED_ONLY_VAL `i_axi_AXI_S7_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S8_ON_AW_SHARED_VAL
  `define AXI_S8_ON_AW_SHARED_VAL `i_axi_AXI_S8_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S8_ON_AW_SHARED_ONLY
  `define AXI_S8_ON_AW_SHARED_ONLY `i_axi_AXI_S8_ON_AW_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S8_ON_AW_SHARED_ONLY_VAL
  `define AXI_S8_ON_AW_SHARED_ONLY_VAL `i_axi_AXI_S8_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S9_ON_AW_SHARED_VAL
  `define AXI_S9_ON_AW_SHARED_VAL `i_axi_AXI_S9_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S9_ON_AW_SHARED_ONLY
  `define AXI_S9_ON_AW_SHARED_ONLY `i_axi_AXI_S9_ON_AW_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S9_ON_AW_SHARED_ONLY_VAL
  `define AXI_S9_ON_AW_SHARED_ONLY_VAL `i_axi_AXI_S9_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S10_ON_AW_SHARED_VAL
  `define AXI_S10_ON_AW_SHARED_VAL `i_axi_AXI_S10_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S10_ON_AW_SHARED_ONLY
  `define AXI_S10_ON_AW_SHARED_ONLY `i_axi_AXI_S10_ON_AW_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S10_ON_AW_SHARED_ONLY_VAL
  `define AXI_S10_ON_AW_SHARED_ONLY_VAL `i_axi_AXI_S10_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S11_ON_AW_SHARED_VAL
  `define AXI_S11_ON_AW_SHARED_VAL `i_axi_AXI_S11_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S11_ON_AW_SHARED_ONLY
  `define AXI_S11_ON_AW_SHARED_ONLY `i_axi_AXI_S11_ON_AW_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S11_ON_AW_SHARED_ONLY_VAL
  `define AXI_S11_ON_AW_SHARED_ONLY_VAL `i_axi_AXI_S11_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S12_ON_AW_SHARED_VAL
  `define AXI_S12_ON_AW_SHARED_VAL `i_axi_AXI_S12_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S12_ON_AW_SHARED_ONLY
  `define AXI_S12_ON_AW_SHARED_ONLY `i_axi_AXI_S12_ON_AW_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S12_ON_AW_SHARED_ONLY_VAL
  `define AXI_S12_ON_AW_SHARED_ONLY_VAL `i_axi_AXI_S12_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S13_ON_AW_SHARED_VAL
  `define AXI_S13_ON_AW_SHARED_VAL `i_axi_AXI_S13_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S13_ON_AW_SHARED_ONLY
  `define AXI_S13_ON_AW_SHARED_ONLY `i_axi_AXI_S13_ON_AW_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S13_ON_AW_SHARED_ONLY_VAL
  `define AXI_S13_ON_AW_SHARED_ONLY_VAL `i_axi_AXI_S13_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S14_ON_AW_SHARED_VAL
  `define AXI_S14_ON_AW_SHARED_VAL `i_axi_AXI_S14_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S14_ON_AW_SHARED_ONLY
  `define AXI_S14_ON_AW_SHARED_ONLY `i_axi_AXI_S14_ON_AW_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S14_ON_AW_SHARED_ONLY_VAL
  `define AXI_S14_ON_AW_SHARED_ONLY_VAL `i_axi_AXI_S14_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S15_ON_AW_SHARED_VAL
  `define AXI_S15_ON_AW_SHARED_VAL `i_axi_AXI_S15_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S15_ON_AW_SHARED_ONLY
  `define AXI_S15_ON_AW_SHARED_ONLY `i_axi_AXI_S15_ON_AW_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S15_ON_AW_SHARED_ONLY_VAL
  `define AXI_S15_ON_AW_SHARED_ONLY_VAL `i_axi_AXI_S15_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S16_ON_AW_SHARED_VAL
  `define AXI_S16_ON_AW_SHARED_VAL `i_axi_AXI_S16_ON_AW_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S16_ON_AW_SHARED_ONLY
  `define AXI_S16_ON_AW_SHARED_ONLY `i_axi_AXI_S16_ON_AW_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S16_ON_AW_SHARED_ONLY_VAL
  `define AXI_S16_ON_AW_SHARED_ONLY_VAL `i_axi_AXI_S16_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M1_ON_W_SHARED_VAL
  `define AXI_M1_ON_W_SHARED_VAL `i_axi_AXI_M1_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M2_ON_W_SHARED_VAL
  `define AXI_M2_ON_W_SHARED_VAL `i_axi_AXI_M2_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M3_ON_W_SHARED_VAL
  `define AXI_M3_ON_W_SHARED_VAL `i_axi_AXI_M3_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M4_ON_W_SHARED_VAL
  `define AXI_M4_ON_W_SHARED_VAL `i_axi_AXI_M4_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M5_ON_W_SHARED_VAL
  `define AXI_M5_ON_W_SHARED_VAL `i_axi_AXI_M5_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M6_ON_W_SHARED_VAL
  `define AXI_M6_ON_W_SHARED_VAL `i_axi_AXI_M6_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M7_ON_W_SHARED_VAL
  `define AXI_M7_ON_W_SHARED_VAL `i_axi_AXI_M7_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M8_ON_W_SHARED_VAL
  `define AXI_M8_ON_W_SHARED_VAL `i_axi_AXI_M8_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M9_ON_W_SHARED_VAL
  `define AXI_M9_ON_W_SHARED_VAL `i_axi_AXI_M9_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M10_ON_W_SHARED_VAL
  `define AXI_M10_ON_W_SHARED_VAL `i_axi_AXI_M10_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M11_ON_W_SHARED_VAL
  `define AXI_M11_ON_W_SHARED_VAL `i_axi_AXI_M11_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M12_ON_W_SHARED_VAL
  `define AXI_M12_ON_W_SHARED_VAL `i_axi_AXI_M12_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M13_ON_W_SHARED_VAL
  `define AXI_M13_ON_W_SHARED_VAL `i_axi_AXI_M13_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M14_ON_W_SHARED_VAL
  `define AXI_M14_ON_W_SHARED_VAL `i_axi_AXI_M14_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M15_ON_W_SHARED_VAL
  `define AXI_M15_ON_W_SHARED_VAL `i_axi_AXI_M15_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M16_ON_W_SHARED_VAL
  `define AXI_M16_ON_W_SHARED_VAL `i_axi_AXI_M16_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S0_ON_W_SHARED_VAL
  `define AXI_S0_ON_W_SHARED_VAL `i_axi_AXI_S0_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S0_ON_W_SHARED_ONLY
  `define AXI_S0_ON_W_SHARED_ONLY `i_axi_AXI_S0_ON_W_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S0_ON_W_SHARED_ONLY_VAL
  `define AXI_S0_ON_W_SHARED_ONLY_VAL `i_axi_AXI_S0_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S1_ON_W_SHARED_VAL
  `define AXI_S1_ON_W_SHARED_VAL `i_axi_AXI_S1_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S1_ON_W_SHARED_ONLY
  `define AXI_S1_ON_W_SHARED_ONLY `i_axi_AXI_S1_ON_W_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S1_ON_W_SHARED_ONLY_VAL
  `define AXI_S1_ON_W_SHARED_ONLY_VAL `i_axi_AXI_S1_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S2_ON_W_SHARED_VAL
  `define AXI_S2_ON_W_SHARED_VAL `i_axi_AXI_S2_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S2_ON_W_SHARED_ONLY
  `define AXI_S2_ON_W_SHARED_ONLY `i_axi_AXI_S2_ON_W_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S2_ON_W_SHARED_ONLY_VAL
  `define AXI_S2_ON_W_SHARED_ONLY_VAL `i_axi_AXI_S2_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S3_ON_W_SHARED_VAL
  `define AXI_S3_ON_W_SHARED_VAL `i_axi_AXI_S3_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S3_ON_W_SHARED_ONLY
  `define AXI_S3_ON_W_SHARED_ONLY `i_axi_AXI_S3_ON_W_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S3_ON_W_SHARED_ONLY_VAL
  `define AXI_S3_ON_W_SHARED_ONLY_VAL `i_axi_AXI_S3_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S4_ON_W_SHARED_VAL
  `define AXI_S4_ON_W_SHARED_VAL `i_axi_AXI_S4_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S4_ON_W_SHARED_ONLY
  `define AXI_S4_ON_W_SHARED_ONLY `i_axi_AXI_S4_ON_W_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S4_ON_W_SHARED_ONLY_VAL
  `define AXI_S4_ON_W_SHARED_ONLY_VAL `i_axi_AXI_S4_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S5_ON_W_SHARED_VAL
  `define AXI_S5_ON_W_SHARED_VAL `i_axi_AXI_S5_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S5_ON_W_SHARED_ONLY
  `define AXI_S5_ON_W_SHARED_ONLY `i_axi_AXI_S5_ON_W_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S5_ON_W_SHARED_ONLY_VAL
  `define AXI_S5_ON_W_SHARED_ONLY_VAL `i_axi_AXI_S5_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S6_ON_W_SHARED_VAL
  `define AXI_S6_ON_W_SHARED_VAL `i_axi_AXI_S6_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S6_ON_W_SHARED_ONLY
  `define AXI_S6_ON_W_SHARED_ONLY `i_axi_AXI_S6_ON_W_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S6_ON_W_SHARED_ONLY_VAL
  `define AXI_S6_ON_W_SHARED_ONLY_VAL `i_axi_AXI_S6_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S7_ON_W_SHARED_VAL
  `define AXI_S7_ON_W_SHARED_VAL `i_axi_AXI_S7_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S7_ON_W_SHARED_ONLY
  `define AXI_S7_ON_W_SHARED_ONLY `i_axi_AXI_S7_ON_W_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S7_ON_W_SHARED_ONLY_VAL
  `define AXI_S7_ON_W_SHARED_ONLY_VAL `i_axi_AXI_S7_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S8_ON_W_SHARED_VAL
  `define AXI_S8_ON_W_SHARED_VAL `i_axi_AXI_S8_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S8_ON_W_SHARED_ONLY
  `define AXI_S8_ON_W_SHARED_ONLY `i_axi_AXI_S8_ON_W_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S8_ON_W_SHARED_ONLY_VAL
  `define AXI_S8_ON_W_SHARED_ONLY_VAL `i_axi_AXI_S8_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S9_ON_W_SHARED_VAL
  `define AXI_S9_ON_W_SHARED_VAL `i_axi_AXI_S9_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S9_ON_W_SHARED_ONLY
  `define AXI_S9_ON_W_SHARED_ONLY `i_axi_AXI_S9_ON_W_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S9_ON_W_SHARED_ONLY_VAL
  `define AXI_S9_ON_W_SHARED_ONLY_VAL `i_axi_AXI_S9_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S10_ON_W_SHARED_VAL
  `define AXI_S10_ON_W_SHARED_VAL `i_axi_AXI_S10_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S10_ON_W_SHARED_ONLY
  `define AXI_S10_ON_W_SHARED_ONLY `i_axi_AXI_S10_ON_W_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S10_ON_W_SHARED_ONLY_VAL
  `define AXI_S10_ON_W_SHARED_ONLY_VAL `i_axi_AXI_S10_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S11_ON_W_SHARED_VAL
  `define AXI_S11_ON_W_SHARED_VAL `i_axi_AXI_S11_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S11_ON_W_SHARED_ONLY
  `define AXI_S11_ON_W_SHARED_ONLY `i_axi_AXI_S11_ON_W_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S11_ON_W_SHARED_ONLY_VAL
  `define AXI_S11_ON_W_SHARED_ONLY_VAL `i_axi_AXI_S11_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S12_ON_W_SHARED_VAL
  `define AXI_S12_ON_W_SHARED_VAL `i_axi_AXI_S12_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S12_ON_W_SHARED_ONLY
  `define AXI_S12_ON_W_SHARED_ONLY `i_axi_AXI_S12_ON_W_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S12_ON_W_SHARED_ONLY_VAL
  `define AXI_S12_ON_W_SHARED_ONLY_VAL `i_axi_AXI_S12_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S13_ON_W_SHARED_VAL
  `define AXI_S13_ON_W_SHARED_VAL `i_axi_AXI_S13_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S13_ON_W_SHARED_ONLY
  `define AXI_S13_ON_W_SHARED_ONLY `i_axi_AXI_S13_ON_W_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S13_ON_W_SHARED_ONLY_VAL
  `define AXI_S13_ON_W_SHARED_ONLY_VAL `i_axi_AXI_S13_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S14_ON_W_SHARED_VAL
  `define AXI_S14_ON_W_SHARED_VAL `i_axi_AXI_S14_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S14_ON_W_SHARED_ONLY
  `define AXI_S14_ON_W_SHARED_ONLY `i_axi_AXI_S14_ON_W_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S14_ON_W_SHARED_ONLY_VAL
  `define AXI_S14_ON_W_SHARED_ONLY_VAL `i_axi_AXI_S14_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S15_ON_W_SHARED_VAL
  `define AXI_S15_ON_W_SHARED_VAL `i_axi_AXI_S15_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S15_ON_W_SHARED_ONLY
  `define AXI_S15_ON_W_SHARED_ONLY `i_axi_AXI_S15_ON_W_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S15_ON_W_SHARED_ONLY_VAL
  `define AXI_S15_ON_W_SHARED_ONLY_VAL `i_axi_AXI_S15_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S16_ON_W_SHARED_VAL
  `define AXI_S16_ON_W_SHARED_VAL `i_axi_AXI_S16_ON_W_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S16_ON_W_SHARED_ONLY
  `define AXI_S16_ON_W_SHARED_ONLY `i_axi_AXI_S16_ON_W_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_S16_ON_W_SHARED_ONLY_VAL
  `define AXI_S16_ON_W_SHARED_ONLY_VAL `i_axi_AXI_S16_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S0_ON_R_SHARED_VAL
  `define AXI_S0_ON_R_SHARED_VAL `i_axi_AXI_S0_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S1_ON_R_SHARED_VAL
  `define AXI_S1_ON_R_SHARED_VAL `i_axi_AXI_S1_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S2_ON_R_SHARED_VAL
  `define AXI_S2_ON_R_SHARED_VAL `i_axi_AXI_S2_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S3_ON_R_SHARED_VAL
  `define AXI_S3_ON_R_SHARED_VAL `i_axi_AXI_S3_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S4_ON_R_SHARED_VAL
  `define AXI_S4_ON_R_SHARED_VAL `i_axi_AXI_S4_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S5_ON_R_SHARED_VAL
  `define AXI_S5_ON_R_SHARED_VAL `i_axi_AXI_S5_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S6_ON_R_SHARED_VAL
  `define AXI_S6_ON_R_SHARED_VAL `i_axi_AXI_S6_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S7_ON_R_SHARED_VAL
  `define AXI_S7_ON_R_SHARED_VAL `i_axi_AXI_S7_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S8_ON_R_SHARED_VAL
  `define AXI_S8_ON_R_SHARED_VAL `i_axi_AXI_S8_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S9_ON_R_SHARED_VAL
  `define AXI_S9_ON_R_SHARED_VAL `i_axi_AXI_S9_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S10_ON_R_SHARED_VAL
  `define AXI_S10_ON_R_SHARED_VAL `i_axi_AXI_S10_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S11_ON_R_SHARED_VAL
  `define AXI_S11_ON_R_SHARED_VAL `i_axi_AXI_S11_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S12_ON_R_SHARED_VAL
  `define AXI_S12_ON_R_SHARED_VAL `i_axi_AXI_S12_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S13_ON_R_SHARED_VAL
  `define AXI_S13_ON_R_SHARED_VAL `i_axi_AXI_S13_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S14_ON_R_SHARED_VAL
  `define AXI_S14_ON_R_SHARED_VAL `i_axi_AXI_S14_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S15_ON_R_SHARED_VAL
  `define AXI_S15_ON_R_SHARED_VAL `i_axi_AXI_S15_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S16_ON_R_SHARED_VAL
  `define AXI_S16_ON_R_SHARED_VAL `i_axi_AXI_S16_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M1_ON_R_SHARED_VAL
  `define AXI_M1_ON_R_SHARED_VAL `i_axi_AXI_M1_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M1_ON_R_SHARED_ONLY
  `define AXI_M1_ON_R_SHARED_ONLY `i_axi_AXI_M1_ON_R_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M1_ON_R_SHARED_ONLY_VAL
  `define AXI_M1_ON_R_SHARED_ONLY_VAL `i_axi_AXI_M1_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M2_ON_R_SHARED_VAL
  `define AXI_M2_ON_R_SHARED_VAL `i_axi_AXI_M2_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M2_ON_R_SHARED_ONLY
  `define AXI_M2_ON_R_SHARED_ONLY `i_axi_AXI_M2_ON_R_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M2_ON_R_SHARED_ONLY_VAL
  `define AXI_M2_ON_R_SHARED_ONLY_VAL `i_axi_AXI_M2_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M3_ON_R_SHARED_VAL
  `define AXI_M3_ON_R_SHARED_VAL `i_axi_AXI_M3_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M3_ON_R_SHARED_ONLY
  `define AXI_M3_ON_R_SHARED_ONLY `i_axi_AXI_M3_ON_R_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M3_ON_R_SHARED_ONLY_VAL
  `define AXI_M3_ON_R_SHARED_ONLY_VAL `i_axi_AXI_M3_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M4_ON_R_SHARED_VAL
  `define AXI_M4_ON_R_SHARED_VAL `i_axi_AXI_M4_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M4_ON_R_SHARED_ONLY
  `define AXI_M4_ON_R_SHARED_ONLY `i_axi_AXI_M4_ON_R_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M4_ON_R_SHARED_ONLY_VAL
  `define AXI_M4_ON_R_SHARED_ONLY_VAL `i_axi_AXI_M4_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M5_ON_R_SHARED_VAL
  `define AXI_M5_ON_R_SHARED_VAL `i_axi_AXI_M5_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M5_ON_R_SHARED_ONLY
  `define AXI_M5_ON_R_SHARED_ONLY `i_axi_AXI_M5_ON_R_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M5_ON_R_SHARED_ONLY_VAL
  `define AXI_M5_ON_R_SHARED_ONLY_VAL `i_axi_AXI_M5_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M6_ON_R_SHARED_VAL
  `define AXI_M6_ON_R_SHARED_VAL `i_axi_AXI_M6_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M6_ON_R_SHARED_ONLY
  `define AXI_M6_ON_R_SHARED_ONLY `i_axi_AXI_M6_ON_R_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M6_ON_R_SHARED_ONLY_VAL
  `define AXI_M6_ON_R_SHARED_ONLY_VAL `i_axi_AXI_M6_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M7_ON_R_SHARED_VAL
  `define AXI_M7_ON_R_SHARED_VAL `i_axi_AXI_M7_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M7_ON_R_SHARED_ONLY
  `define AXI_M7_ON_R_SHARED_ONLY `i_axi_AXI_M7_ON_R_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M7_ON_R_SHARED_ONLY_VAL
  `define AXI_M7_ON_R_SHARED_ONLY_VAL `i_axi_AXI_M7_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M8_ON_R_SHARED_VAL
  `define AXI_M8_ON_R_SHARED_VAL `i_axi_AXI_M8_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M8_ON_R_SHARED_ONLY
  `define AXI_M8_ON_R_SHARED_ONLY `i_axi_AXI_M8_ON_R_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M8_ON_R_SHARED_ONLY_VAL
  `define AXI_M8_ON_R_SHARED_ONLY_VAL `i_axi_AXI_M8_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M9_ON_R_SHARED_VAL
  `define AXI_M9_ON_R_SHARED_VAL `i_axi_AXI_M9_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M9_ON_R_SHARED_ONLY
  `define AXI_M9_ON_R_SHARED_ONLY `i_axi_AXI_M9_ON_R_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M9_ON_R_SHARED_ONLY_VAL
  `define AXI_M9_ON_R_SHARED_ONLY_VAL `i_axi_AXI_M9_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M10_ON_R_SHARED_VAL
  `define AXI_M10_ON_R_SHARED_VAL `i_axi_AXI_M10_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M10_ON_R_SHARED_ONLY
  `define AXI_M10_ON_R_SHARED_ONLY `i_axi_AXI_M10_ON_R_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M10_ON_R_SHARED_ONLY_VAL
  `define AXI_M10_ON_R_SHARED_ONLY_VAL `i_axi_AXI_M10_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M11_ON_R_SHARED_VAL
  `define AXI_M11_ON_R_SHARED_VAL `i_axi_AXI_M11_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M11_ON_R_SHARED_ONLY
  `define AXI_M11_ON_R_SHARED_ONLY `i_axi_AXI_M11_ON_R_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M11_ON_R_SHARED_ONLY_VAL
  `define AXI_M11_ON_R_SHARED_ONLY_VAL `i_axi_AXI_M11_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M12_ON_R_SHARED_VAL
  `define AXI_M12_ON_R_SHARED_VAL `i_axi_AXI_M12_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M12_ON_R_SHARED_ONLY
  `define AXI_M12_ON_R_SHARED_ONLY `i_axi_AXI_M12_ON_R_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M12_ON_R_SHARED_ONLY_VAL
  `define AXI_M12_ON_R_SHARED_ONLY_VAL `i_axi_AXI_M12_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M13_ON_R_SHARED_VAL
  `define AXI_M13_ON_R_SHARED_VAL `i_axi_AXI_M13_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M13_ON_R_SHARED_ONLY
  `define AXI_M13_ON_R_SHARED_ONLY `i_axi_AXI_M13_ON_R_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M13_ON_R_SHARED_ONLY_VAL
  `define AXI_M13_ON_R_SHARED_ONLY_VAL `i_axi_AXI_M13_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M14_ON_R_SHARED_VAL
  `define AXI_M14_ON_R_SHARED_VAL `i_axi_AXI_M14_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M14_ON_R_SHARED_ONLY
  `define AXI_M14_ON_R_SHARED_ONLY `i_axi_AXI_M14_ON_R_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M14_ON_R_SHARED_ONLY_VAL
  `define AXI_M14_ON_R_SHARED_ONLY_VAL `i_axi_AXI_M14_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M15_ON_R_SHARED_VAL
  `define AXI_M15_ON_R_SHARED_VAL `i_axi_AXI_M15_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M15_ON_R_SHARED_ONLY
  `define AXI_M15_ON_R_SHARED_ONLY `i_axi_AXI_M15_ON_R_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M15_ON_R_SHARED_ONLY_VAL
  `define AXI_M15_ON_R_SHARED_ONLY_VAL `i_axi_AXI_M15_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M16_ON_R_SHARED_VAL
  `define AXI_M16_ON_R_SHARED_VAL `i_axi_AXI_M16_ON_R_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M16_ON_R_SHARED_ONLY
  `define AXI_M16_ON_R_SHARED_ONLY `i_axi_AXI_M16_ON_R_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M16_ON_R_SHARED_ONLY_VAL
  `define AXI_M16_ON_R_SHARED_ONLY_VAL `i_axi_AXI_M16_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_S0_ON_B_SHARED_VAL
  `define AXI_S0_ON_B_SHARED_VAL `i_axi_AXI_S0_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S1_ON_B_SHARED_VAL
  `define AXI_S1_ON_B_SHARED_VAL `i_axi_AXI_S1_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S2_ON_B_SHARED_VAL
  `define AXI_S2_ON_B_SHARED_VAL `i_axi_AXI_S2_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S3_ON_B_SHARED_VAL
  `define AXI_S3_ON_B_SHARED_VAL `i_axi_AXI_S3_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S4_ON_B_SHARED_VAL
  `define AXI_S4_ON_B_SHARED_VAL `i_axi_AXI_S4_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S5_ON_B_SHARED_VAL
  `define AXI_S5_ON_B_SHARED_VAL `i_axi_AXI_S5_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S6_ON_B_SHARED_VAL
  `define AXI_S6_ON_B_SHARED_VAL `i_axi_AXI_S6_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S7_ON_B_SHARED_VAL
  `define AXI_S7_ON_B_SHARED_VAL `i_axi_AXI_S7_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S8_ON_B_SHARED_VAL
  `define AXI_S8_ON_B_SHARED_VAL `i_axi_AXI_S8_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S9_ON_B_SHARED_VAL
  `define AXI_S9_ON_B_SHARED_VAL `i_axi_AXI_S9_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S10_ON_B_SHARED_VAL
  `define AXI_S10_ON_B_SHARED_VAL `i_axi_AXI_S10_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S11_ON_B_SHARED_VAL
  `define AXI_S11_ON_B_SHARED_VAL `i_axi_AXI_S11_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S12_ON_B_SHARED_VAL
  `define AXI_S12_ON_B_SHARED_VAL `i_axi_AXI_S12_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S13_ON_B_SHARED_VAL
  `define AXI_S13_ON_B_SHARED_VAL `i_axi_AXI_S13_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S14_ON_B_SHARED_VAL
  `define AXI_S14_ON_B_SHARED_VAL `i_axi_AXI_S14_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S15_ON_B_SHARED_VAL
  `define AXI_S15_ON_B_SHARED_VAL `i_axi_AXI_S15_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_S16_ON_B_SHARED_VAL
  `define AXI_S16_ON_B_SHARED_VAL `i_axi_AXI_S16_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M1_ON_B_SHARED_VAL
  `define AXI_M1_ON_B_SHARED_VAL `i_axi_AXI_M1_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M1_ON_B_SHARED_ONLY
  `define AXI_M1_ON_B_SHARED_ONLY `i_axi_AXI_M1_ON_B_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M1_ON_B_SHARED_ONLY_VAL
  `define AXI_M1_ON_B_SHARED_ONLY_VAL `i_axi_AXI_M1_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M2_ON_B_SHARED_VAL
  `define AXI_M2_ON_B_SHARED_VAL `i_axi_AXI_M2_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M2_ON_B_SHARED_ONLY
  `define AXI_M2_ON_B_SHARED_ONLY `i_axi_AXI_M2_ON_B_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M2_ON_B_SHARED_ONLY_VAL
  `define AXI_M2_ON_B_SHARED_ONLY_VAL `i_axi_AXI_M2_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M3_ON_B_SHARED_VAL
  `define AXI_M3_ON_B_SHARED_VAL `i_axi_AXI_M3_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M3_ON_B_SHARED_ONLY
  `define AXI_M3_ON_B_SHARED_ONLY `i_axi_AXI_M3_ON_B_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M3_ON_B_SHARED_ONLY_VAL
  `define AXI_M3_ON_B_SHARED_ONLY_VAL `i_axi_AXI_M3_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M4_ON_B_SHARED_VAL
  `define AXI_M4_ON_B_SHARED_VAL `i_axi_AXI_M4_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M4_ON_B_SHARED_ONLY
  `define AXI_M4_ON_B_SHARED_ONLY `i_axi_AXI_M4_ON_B_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M4_ON_B_SHARED_ONLY_VAL
  `define AXI_M4_ON_B_SHARED_ONLY_VAL `i_axi_AXI_M4_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M5_ON_B_SHARED_VAL
  `define AXI_M5_ON_B_SHARED_VAL `i_axi_AXI_M5_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M5_ON_B_SHARED_ONLY
  `define AXI_M5_ON_B_SHARED_ONLY `i_axi_AXI_M5_ON_B_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M5_ON_B_SHARED_ONLY_VAL
  `define AXI_M5_ON_B_SHARED_ONLY_VAL `i_axi_AXI_M5_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M6_ON_B_SHARED_VAL
  `define AXI_M6_ON_B_SHARED_VAL `i_axi_AXI_M6_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M6_ON_B_SHARED_ONLY
  `define AXI_M6_ON_B_SHARED_ONLY `i_axi_AXI_M6_ON_B_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M6_ON_B_SHARED_ONLY_VAL
  `define AXI_M6_ON_B_SHARED_ONLY_VAL `i_axi_AXI_M6_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M7_ON_B_SHARED_VAL
  `define AXI_M7_ON_B_SHARED_VAL `i_axi_AXI_M7_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M7_ON_B_SHARED_ONLY
  `define AXI_M7_ON_B_SHARED_ONLY `i_axi_AXI_M7_ON_B_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M7_ON_B_SHARED_ONLY_VAL
  `define AXI_M7_ON_B_SHARED_ONLY_VAL `i_axi_AXI_M7_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M8_ON_B_SHARED_VAL
  `define AXI_M8_ON_B_SHARED_VAL `i_axi_AXI_M8_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M8_ON_B_SHARED_ONLY
  `define AXI_M8_ON_B_SHARED_ONLY `i_axi_AXI_M8_ON_B_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M8_ON_B_SHARED_ONLY_VAL
  `define AXI_M8_ON_B_SHARED_ONLY_VAL `i_axi_AXI_M8_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M9_ON_B_SHARED_VAL
  `define AXI_M9_ON_B_SHARED_VAL `i_axi_AXI_M9_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M9_ON_B_SHARED_ONLY
  `define AXI_M9_ON_B_SHARED_ONLY `i_axi_AXI_M9_ON_B_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M9_ON_B_SHARED_ONLY_VAL
  `define AXI_M9_ON_B_SHARED_ONLY_VAL `i_axi_AXI_M9_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M10_ON_B_SHARED_VAL
  `define AXI_M10_ON_B_SHARED_VAL `i_axi_AXI_M10_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M10_ON_B_SHARED_ONLY
  `define AXI_M10_ON_B_SHARED_ONLY `i_axi_AXI_M10_ON_B_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M10_ON_B_SHARED_ONLY_VAL
  `define AXI_M10_ON_B_SHARED_ONLY_VAL `i_axi_AXI_M10_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M11_ON_B_SHARED_VAL
  `define AXI_M11_ON_B_SHARED_VAL `i_axi_AXI_M11_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M11_ON_B_SHARED_ONLY
  `define AXI_M11_ON_B_SHARED_ONLY `i_axi_AXI_M11_ON_B_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M11_ON_B_SHARED_ONLY_VAL
  `define AXI_M11_ON_B_SHARED_ONLY_VAL `i_axi_AXI_M11_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M12_ON_B_SHARED_VAL
  `define AXI_M12_ON_B_SHARED_VAL `i_axi_AXI_M12_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M12_ON_B_SHARED_ONLY
  `define AXI_M12_ON_B_SHARED_ONLY `i_axi_AXI_M12_ON_B_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M12_ON_B_SHARED_ONLY_VAL
  `define AXI_M12_ON_B_SHARED_ONLY_VAL `i_axi_AXI_M12_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M13_ON_B_SHARED_VAL
  `define AXI_M13_ON_B_SHARED_VAL `i_axi_AXI_M13_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M13_ON_B_SHARED_ONLY
  `define AXI_M13_ON_B_SHARED_ONLY `i_axi_AXI_M13_ON_B_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M13_ON_B_SHARED_ONLY_VAL
  `define AXI_M13_ON_B_SHARED_ONLY_VAL `i_axi_AXI_M13_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M14_ON_B_SHARED_VAL
  `define AXI_M14_ON_B_SHARED_VAL `i_axi_AXI_M14_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M14_ON_B_SHARED_ONLY
  `define AXI_M14_ON_B_SHARED_ONLY `i_axi_AXI_M14_ON_B_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M14_ON_B_SHARED_ONLY_VAL
  `define AXI_M14_ON_B_SHARED_ONLY_VAL `i_axi_AXI_M14_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M15_ON_B_SHARED_VAL
  `define AXI_M15_ON_B_SHARED_VAL `i_axi_AXI_M15_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M15_ON_B_SHARED_ONLY
  `define AXI_M15_ON_B_SHARED_ONLY `i_axi_AXI_M15_ON_B_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M15_ON_B_SHARED_ONLY_VAL
  `define AXI_M15_ON_B_SHARED_ONLY_VAL `i_axi_AXI_M15_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_M16_ON_B_SHARED_VAL
  `define AXI_M16_ON_B_SHARED_VAL `i_axi_AXI_M16_ON_B_SHARED_VAL
`endif 

`ifdef i_axi_AXI_M16_ON_B_SHARED_ONLY
  `define AXI_M16_ON_B_SHARED_ONLY `i_axi_AXI_M16_ON_B_SHARED_ONLY
`endif 

`ifdef i_axi_AXI_M16_ON_B_SHARED_ONLY_VAL
  `define AXI_M16_ON_B_SHARED_ONLY_VAL `i_axi_AXI_M16_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef i_axi_AXI_AW_SHARED_PL
  `define AXI_AW_SHARED_PL `i_axi_AXI_AW_SHARED_PL
`endif 

`ifdef i_axi_AXI_AR_SHARED_PL
  `define AXI_AR_SHARED_PL `i_axi_AXI_AR_SHARED_PL
`endif 

`ifdef i_axi_AXI_W_SHARED_PL
  `define AXI_W_SHARED_PL `i_axi_AXI_W_SHARED_PL
`endif 

`ifdef i_axi_AXI_R_SHARED_PL
  `define AXI_R_SHARED_PL `i_axi_AXI_R_SHARED_PL
`endif 

`ifdef i_axi_AXI_B_SHARED_PL
  `define AXI_B_SHARED_PL `i_axi_AXI_B_SHARED_PL
`endif 

`ifdef i_axi_AXI_MCA_HLD_PRIOR
  `define AXI_MCA_HLD_PRIOR `i_axi_AXI_MCA_HLD_PRIOR
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_S0
  `define AXI_AR_MCA_NC_S0 `i_axi_AXI_AR_MCA_NC_S0
`endif 

`ifdef i_axi_AXI_AR_MCA_EN_S0
  `define AXI_AR_MCA_EN_S0 `i_axi_AXI_AR_MCA_EN_S0
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_W_S0
  `define AXI_AR_MCA_NC_W_S0 `i_axi_AXI_AR_MCA_NC_W_S0
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_S0
  `define AXI_AW_MCA_NC_S0 `i_axi_AXI_AW_MCA_NC_S0
`endif 

`ifdef i_axi_AXI_AW_MCA_EN_S0
  `define AXI_AW_MCA_EN_S0 `i_axi_AXI_AW_MCA_EN_S0
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_W_S0
  `define AXI_AW_MCA_NC_W_S0 `i_axi_AXI_AW_MCA_NC_W_S0
`endif 

`ifdef i_axi_AXI_W_MCA_NC_S0
  `define AXI_W_MCA_NC_S0 `i_axi_AXI_W_MCA_NC_S0
`endif 

`ifdef i_axi_AXI_W_MCA_EN_S0
  `define AXI_W_MCA_EN_S0 `i_axi_AXI_W_MCA_EN_S0
`endif 

`ifdef i_axi_AXI_W_MCA_NC_W_S0
  `define AXI_W_MCA_NC_W_S0 `i_axi_AXI_W_MCA_NC_W_S0
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_S1
  `define AXI_AR_MCA_NC_S1 `i_axi_AXI_AR_MCA_NC_S1
`endif 

`ifdef i_axi_AXI_AR_MCA_EN_S1
  `define AXI_AR_MCA_EN_S1 `i_axi_AXI_AR_MCA_EN_S1
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_W_S1
  `define AXI_AR_MCA_NC_W_S1 `i_axi_AXI_AR_MCA_NC_W_S1
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_S1
  `define AXI_AW_MCA_NC_S1 `i_axi_AXI_AW_MCA_NC_S1
`endif 

`ifdef i_axi_AXI_AW_MCA_EN_S1
  `define AXI_AW_MCA_EN_S1 `i_axi_AXI_AW_MCA_EN_S1
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_W_S1
  `define AXI_AW_MCA_NC_W_S1 `i_axi_AXI_AW_MCA_NC_W_S1
`endif 

`ifdef i_axi_AXI_W_MCA_NC_S1
  `define AXI_W_MCA_NC_S1 `i_axi_AXI_W_MCA_NC_S1
`endif 

`ifdef i_axi_AXI_W_MCA_EN_S1
  `define AXI_W_MCA_EN_S1 `i_axi_AXI_W_MCA_EN_S1
`endif 

`ifdef i_axi_AXI_W_MCA_NC_W_S1
  `define AXI_W_MCA_NC_W_S1 `i_axi_AXI_W_MCA_NC_W_S1
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_S2
  `define AXI_AR_MCA_NC_S2 `i_axi_AXI_AR_MCA_NC_S2
`endif 

`ifdef i_axi_AXI_AR_MCA_EN_S2
  `define AXI_AR_MCA_EN_S2 `i_axi_AXI_AR_MCA_EN_S2
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_W_S2
  `define AXI_AR_MCA_NC_W_S2 `i_axi_AXI_AR_MCA_NC_W_S2
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_S2
  `define AXI_AW_MCA_NC_S2 `i_axi_AXI_AW_MCA_NC_S2
`endif 

`ifdef i_axi_AXI_AW_MCA_EN_S2
  `define AXI_AW_MCA_EN_S2 `i_axi_AXI_AW_MCA_EN_S2
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_W_S2
  `define AXI_AW_MCA_NC_W_S2 `i_axi_AXI_AW_MCA_NC_W_S2
`endif 

`ifdef i_axi_AXI_W_MCA_NC_S2
  `define AXI_W_MCA_NC_S2 `i_axi_AXI_W_MCA_NC_S2
`endif 

`ifdef i_axi_AXI_W_MCA_EN_S2
  `define AXI_W_MCA_EN_S2 `i_axi_AXI_W_MCA_EN_S2
`endif 

`ifdef i_axi_AXI_W_MCA_NC_W_S2
  `define AXI_W_MCA_NC_W_S2 `i_axi_AXI_W_MCA_NC_W_S2
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_S3
  `define AXI_AR_MCA_NC_S3 `i_axi_AXI_AR_MCA_NC_S3
`endif 

`ifdef i_axi_AXI_AR_MCA_EN_S3
  `define AXI_AR_MCA_EN_S3 `i_axi_AXI_AR_MCA_EN_S3
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_W_S3
  `define AXI_AR_MCA_NC_W_S3 `i_axi_AXI_AR_MCA_NC_W_S3
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_S3
  `define AXI_AW_MCA_NC_S3 `i_axi_AXI_AW_MCA_NC_S3
`endif 

`ifdef i_axi_AXI_AW_MCA_EN_S3
  `define AXI_AW_MCA_EN_S3 `i_axi_AXI_AW_MCA_EN_S3
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_W_S3
  `define AXI_AW_MCA_NC_W_S3 `i_axi_AXI_AW_MCA_NC_W_S3
`endif 

`ifdef i_axi_AXI_W_MCA_NC_S3
  `define AXI_W_MCA_NC_S3 `i_axi_AXI_W_MCA_NC_S3
`endif 

`ifdef i_axi_AXI_W_MCA_EN_S3
  `define AXI_W_MCA_EN_S3 `i_axi_AXI_W_MCA_EN_S3
`endif 

`ifdef i_axi_AXI_W_MCA_NC_W_S3
  `define AXI_W_MCA_NC_W_S3 `i_axi_AXI_W_MCA_NC_W_S3
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_S4
  `define AXI_AR_MCA_NC_S4 `i_axi_AXI_AR_MCA_NC_S4
`endif 

`ifdef i_axi_AXI_AR_MCA_EN_S4
  `define AXI_AR_MCA_EN_S4 `i_axi_AXI_AR_MCA_EN_S4
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_W_S4
  `define AXI_AR_MCA_NC_W_S4 `i_axi_AXI_AR_MCA_NC_W_S4
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_S4
  `define AXI_AW_MCA_NC_S4 `i_axi_AXI_AW_MCA_NC_S4
`endif 

`ifdef i_axi_AXI_AW_MCA_EN_S4
  `define AXI_AW_MCA_EN_S4 `i_axi_AXI_AW_MCA_EN_S4
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_W_S4
  `define AXI_AW_MCA_NC_W_S4 `i_axi_AXI_AW_MCA_NC_W_S4
`endif 

`ifdef i_axi_AXI_W_MCA_NC_S4
  `define AXI_W_MCA_NC_S4 `i_axi_AXI_W_MCA_NC_S4
`endif 

`ifdef i_axi_AXI_W_MCA_EN_S4
  `define AXI_W_MCA_EN_S4 `i_axi_AXI_W_MCA_EN_S4
`endif 

`ifdef i_axi_AXI_W_MCA_NC_W_S4
  `define AXI_W_MCA_NC_W_S4 `i_axi_AXI_W_MCA_NC_W_S4
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_S5
  `define AXI_AR_MCA_NC_S5 `i_axi_AXI_AR_MCA_NC_S5
`endif 

`ifdef i_axi_AXI_AR_MCA_EN_S5
  `define AXI_AR_MCA_EN_S5 `i_axi_AXI_AR_MCA_EN_S5
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_W_S5
  `define AXI_AR_MCA_NC_W_S5 `i_axi_AXI_AR_MCA_NC_W_S5
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_S5
  `define AXI_AW_MCA_NC_S5 `i_axi_AXI_AW_MCA_NC_S5
`endif 

`ifdef i_axi_AXI_AW_MCA_EN_S5
  `define AXI_AW_MCA_EN_S5 `i_axi_AXI_AW_MCA_EN_S5
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_W_S5
  `define AXI_AW_MCA_NC_W_S5 `i_axi_AXI_AW_MCA_NC_W_S5
`endif 

`ifdef i_axi_AXI_W_MCA_NC_S5
  `define AXI_W_MCA_NC_S5 `i_axi_AXI_W_MCA_NC_S5
`endif 

`ifdef i_axi_AXI_W_MCA_EN_S5
  `define AXI_W_MCA_EN_S5 `i_axi_AXI_W_MCA_EN_S5
`endif 

`ifdef i_axi_AXI_W_MCA_NC_W_S5
  `define AXI_W_MCA_NC_W_S5 `i_axi_AXI_W_MCA_NC_W_S5
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_S6
  `define AXI_AR_MCA_NC_S6 `i_axi_AXI_AR_MCA_NC_S6
`endif 

`ifdef i_axi_AXI_AR_MCA_EN_S6
  `define AXI_AR_MCA_EN_S6 `i_axi_AXI_AR_MCA_EN_S6
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_W_S6
  `define AXI_AR_MCA_NC_W_S6 `i_axi_AXI_AR_MCA_NC_W_S6
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_S6
  `define AXI_AW_MCA_NC_S6 `i_axi_AXI_AW_MCA_NC_S6
`endif 

`ifdef i_axi_AXI_AW_MCA_EN_S6
  `define AXI_AW_MCA_EN_S6 `i_axi_AXI_AW_MCA_EN_S6
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_W_S6
  `define AXI_AW_MCA_NC_W_S6 `i_axi_AXI_AW_MCA_NC_W_S6
`endif 

`ifdef i_axi_AXI_W_MCA_NC_S6
  `define AXI_W_MCA_NC_S6 `i_axi_AXI_W_MCA_NC_S6
`endif 

`ifdef i_axi_AXI_W_MCA_EN_S6
  `define AXI_W_MCA_EN_S6 `i_axi_AXI_W_MCA_EN_S6
`endif 

`ifdef i_axi_AXI_W_MCA_NC_W_S6
  `define AXI_W_MCA_NC_W_S6 `i_axi_AXI_W_MCA_NC_W_S6
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_S7
  `define AXI_AR_MCA_NC_S7 `i_axi_AXI_AR_MCA_NC_S7
`endif 

`ifdef i_axi_AXI_AR_MCA_EN_S7
  `define AXI_AR_MCA_EN_S7 `i_axi_AXI_AR_MCA_EN_S7
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_W_S7
  `define AXI_AR_MCA_NC_W_S7 `i_axi_AXI_AR_MCA_NC_W_S7
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_S7
  `define AXI_AW_MCA_NC_S7 `i_axi_AXI_AW_MCA_NC_S7
`endif 

`ifdef i_axi_AXI_AW_MCA_EN_S7
  `define AXI_AW_MCA_EN_S7 `i_axi_AXI_AW_MCA_EN_S7
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_W_S7
  `define AXI_AW_MCA_NC_W_S7 `i_axi_AXI_AW_MCA_NC_W_S7
`endif 

`ifdef i_axi_AXI_W_MCA_NC_S7
  `define AXI_W_MCA_NC_S7 `i_axi_AXI_W_MCA_NC_S7
`endif 

`ifdef i_axi_AXI_W_MCA_EN_S7
  `define AXI_W_MCA_EN_S7 `i_axi_AXI_W_MCA_EN_S7
`endif 

`ifdef i_axi_AXI_W_MCA_NC_W_S7
  `define AXI_W_MCA_NC_W_S7 `i_axi_AXI_W_MCA_NC_W_S7
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_S8
  `define AXI_AR_MCA_NC_S8 `i_axi_AXI_AR_MCA_NC_S8
`endif 

`ifdef i_axi_AXI_AR_MCA_EN_S8
  `define AXI_AR_MCA_EN_S8 `i_axi_AXI_AR_MCA_EN_S8
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_W_S8
  `define AXI_AR_MCA_NC_W_S8 `i_axi_AXI_AR_MCA_NC_W_S8
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_S8
  `define AXI_AW_MCA_NC_S8 `i_axi_AXI_AW_MCA_NC_S8
`endif 

`ifdef i_axi_AXI_AW_MCA_EN_S8
  `define AXI_AW_MCA_EN_S8 `i_axi_AXI_AW_MCA_EN_S8
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_W_S8
  `define AXI_AW_MCA_NC_W_S8 `i_axi_AXI_AW_MCA_NC_W_S8
`endif 

`ifdef i_axi_AXI_W_MCA_NC_S8
  `define AXI_W_MCA_NC_S8 `i_axi_AXI_W_MCA_NC_S8
`endif 

`ifdef i_axi_AXI_W_MCA_EN_S8
  `define AXI_W_MCA_EN_S8 `i_axi_AXI_W_MCA_EN_S8
`endif 

`ifdef i_axi_AXI_W_MCA_NC_W_S8
  `define AXI_W_MCA_NC_W_S8 `i_axi_AXI_W_MCA_NC_W_S8
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_S9
  `define AXI_AR_MCA_NC_S9 `i_axi_AXI_AR_MCA_NC_S9
`endif 

`ifdef i_axi_AXI_AR_MCA_EN_S9
  `define AXI_AR_MCA_EN_S9 `i_axi_AXI_AR_MCA_EN_S9
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_W_S9
  `define AXI_AR_MCA_NC_W_S9 `i_axi_AXI_AR_MCA_NC_W_S9
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_S9
  `define AXI_AW_MCA_NC_S9 `i_axi_AXI_AW_MCA_NC_S9
`endif 

`ifdef i_axi_AXI_AW_MCA_EN_S9
  `define AXI_AW_MCA_EN_S9 `i_axi_AXI_AW_MCA_EN_S9
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_W_S9
  `define AXI_AW_MCA_NC_W_S9 `i_axi_AXI_AW_MCA_NC_W_S9
`endif 

`ifdef i_axi_AXI_W_MCA_NC_S9
  `define AXI_W_MCA_NC_S9 `i_axi_AXI_W_MCA_NC_S9
`endif 

`ifdef i_axi_AXI_W_MCA_EN_S9
  `define AXI_W_MCA_EN_S9 `i_axi_AXI_W_MCA_EN_S9
`endif 

`ifdef i_axi_AXI_W_MCA_NC_W_S9
  `define AXI_W_MCA_NC_W_S9 `i_axi_AXI_W_MCA_NC_W_S9
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_S10
  `define AXI_AR_MCA_NC_S10 `i_axi_AXI_AR_MCA_NC_S10
`endif 

`ifdef i_axi_AXI_AR_MCA_EN_S10
  `define AXI_AR_MCA_EN_S10 `i_axi_AXI_AR_MCA_EN_S10
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_W_S10
  `define AXI_AR_MCA_NC_W_S10 `i_axi_AXI_AR_MCA_NC_W_S10
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_S10
  `define AXI_AW_MCA_NC_S10 `i_axi_AXI_AW_MCA_NC_S10
`endif 

`ifdef i_axi_AXI_AW_MCA_EN_S10
  `define AXI_AW_MCA_EN_S10 `i_axi_AXI_AW_MCA_EN_S10
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_W_S10
  `define AXI_AW_MCA_NC_W_S10 `i_axi_AXI_AW_MCA_NC_W_S10
`endif 

`ifdef i_axi_AXI_W_MCA_NC_S10
  `define AXI_W_MCA_NC_S10 `i_axi_AXI_W_MCA_NC_S10
`endif 

`ifdef i_axi_AXI_W_MCA_EN_S10
  `define AXI_W_MCA_EN_S10 `i_axi_AXI_W_MCA_EN_S10
`endif 

`ifdef i_axi_AXI_W_MCA_NC_W_S10
  `define AXI_W_MCA_NC_W_S10 `i_axi_AXI_W_MCA_NC_W_S10
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_S11
  `define AXI_AR_MCA_NC_S11 `i_axi_AXI_AR_MCA_NC_S11
`endif 

`ifdef i_axi_AXI_AR_MCA_EN_S11
  `define AXI_AR_MCA_EN_S11 `i_axi_AXI_AR_MCA_EN_S11
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_W_S11
  `define AXI_AR_MCA_NC_W_S11 `i_axi_AXI_AR_MCA_NC_W_S11
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_S11
  `define AXI_AW_MCA_NC_S11 `i_axi_AXI_AW_MCA_NC_S11
`endif 

`ifdef i_axi_AXI_AW_MCA_EN_S11
  `define AXI_AW_MCA_EN_S11 `i_axi_AXI_AW_MCA_EN_S11
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_W_S11
  `define AXI_AW_MCA_NC_W_S11 `i_axi_AXI_AW_MCA_NC_W_S11
`endif 

`ifdef i_axi_AXI_W_MCA_NC_S11
  `define AXI_W_MCA_NC_S11 `i_axi_AXI_W_MCA_NC_S11
`endif 

`ifdef i_axi_AXI_W_MCA_EN_S11
  `define AXI_W_MCA_EN_S11 `i_axi_AXI_W_MCA_EN_S11
`endif 

`ifdef i_axi_AXI_W_MCA_NC_W_S11
  `define AXI_W_MCA_NC_W_S11 `i_axi_AXI_W_MCA_NC_W_S11
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_S12
  `define AXI_AR_MCA_NC_S12 `i_axi_AXI_AR_MCA_NC_S12
`endif 

`ifdef i_axi_AXI_AR_MCA_EN_S12
  `define AXI_AR_MCA_EN_S12 `i_axi_AXI_AR_MCA_EN_S12
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_W_S12
  `define AXI_AR_MCA_NC_W_S12 `i_axi_AXI_AR_MCA_NC_W_S12
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_S12
  `define AXI_AW_MCA_NC_S12 `i_axi_AXI_AW_MCA_NC_S12
`endif 

`ifdef i_axi_AXI_AW_MCA_EN_S12
  `define AXI_AW_MCA_EN_S12 `i_axi_AXI_AW_MCA_EN_S12
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_W_S12
  `define AXI_AW_MCA_NC_W_S12 `i_axi_AXI_AW_MCA_NC_W_S12
`endif 

`ifdef i_axi_AXI_W_MCA_NC_S12
  `define AXI_W_MCA_NC_S12 `i_axi_AXI_W_MCA_NC_S12
`endif 

`ifdef i_axi_AXI_W_MCA_EN_S12
  `define AXI_W_MCA_EN_S12 `i_axi_AXI_W_MCA_EN_S12
`endif 

`ifdef i_axi_AXI_W_MCA_NC_W_S12
  `define AXI_W_MCA_NC_W_S12 `i_axi_AXI_W_MCA_NC_W_S12
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_S13
  `define AXI_AR_MCA_NC_S13 `i_axi_AXI_AR_MCA_NC_S13
`endif 

`ifdef i_axi_AXI_AR_MCA_EN_S13
  `define AXI_AR_MCA_EN_S13 `i_axi_AXI_AR_MCA_EN_S13
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_W_S13
  `define AXI_AR_MCA_NC_W_S13 `i_axi_AXI_AR_MCA_NC_W_S13
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_S13
  `define AXI_AW_MCA_NC_S13 `i_axi_AXI_AW_MCA_NC_S13
`endif 

`ifdef i_axi_AXI_AW_MCA_EN_S13
  `define AXI_AW_MCA_EN_S13 `i_axi_AXI_AW_MCA_EN_S13
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_W_S13
  `define AXI_AW_MCA_NC_W_S13 `i_axi_AXI_AW_MCA_NC_W_S13
`endif 

`ifdef i_axi_AXI_W_MCA_NC_S13
  `define AXI_W_MCA_NC_S13 `i_axi_AXI_W_MCA_NC_S13
`endif 

`ifdef i_axi_AXI_W_MCA_EN_S13
  `define AXI_W_MCA_EN_S13 `i_axi_AXI_W_MCA_EN_S13
`endif 

`ifdef i_axi_AXI_W_MCA_NC_W_S13
  `define AXI_W_MCA_NC_W_S13 `i_axi_AXI_W_MCA_NC_W_S13
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_S14
  `define AXI_AR_MCA_NC_S14 `i_axi_AXI_AR_MCA_NC_S14
`endif 

`ifdef i_axi_AXI_AR_MCA_EN_S14
  `define AXI_AR_MCA_EN_S14 `i_axi_AXI_AR_MCA_EN_S14
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_W_S14
  `define AXI_AR_MCA_NC_W_S14 `i_axi_AXI_AR_MCA_NC_W_S14
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_S14
  `define AXI_AW_MCA_NC_S14 `i_axi_AXI_AW_MCA_NC_S14
`endif 

`ifdef i_axi_AXI_AW_MCA_EN_S14
  `define AXI_AW_MCA_EN_S14 `i_axi_AXI_AW_MCA_EN_S14
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_W_S14
  `define AXI_AW_MCA_NC_W_S14 `i_axi_AXI_AW_MCA_NC_W_S14
`endif 

`ifdef i_axi_AXI_W_MCA_NC_S14
  `define AXI_W_MCA_NC_S14 `i_axi_AXI_W_MCA_NC_S14
`endif 

`ifdef i_axi_AXI_W_MCA_EN_S14
  `define AXI_W_MCA_EN_S14 `i_axi_AXI_W_MCA_EN_S14
`endif 

`ifdef i_axi_AXI_W_MCA_NC_W_S14
  `define AXI_W_MCA_NC_W_S14 `i_axi_AXI_W_MCA_NC_W_S14
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_S15
  `define AXI_AR_MCA_NC_S15 `i_axi_AXI_AR_MCA_NC_S15
`endif 

`ifdef i_axi_AXI_AR_MCA_EN_S15
  `define AXI_AR_MCA_EN_S15 `i_axi_AXI_AR_MCA_EN_S15
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_W_S15
  `define AXI_AR_MCA_NC_W_S15 `i_axi_AXI_AR_MCA_NC_W_S15
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_S15
  `define AXI_AW_MCA_NC_S15 `i_axi_AXI_AW_MCA_NC_S15
`endif 

`ifdef i_axi_AXI_AW_MCA_EN_S15
  `define AXI_AW_MCA_EN_S15 `i_axi_AXI_AW_MCA_EN_S15
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_W_S15
  `define AXI_AW_MCA_NC_W_S15 `i_axi_AXI_AW_MCA_NC_W_S15
`endif 

`ifdef i_axi_AXI_W_MCA_NC_S15
  `define AXI_W_MCA_NC_S15 `i_axi_AXI_W_MCA_NC_S15
`endif 

`ifdef i_axi_AXI_W_MCA_EN_S15
  `define AXI_W_MCA_EN_S15 `i_axi_AXI_W_MCA_EN_S15
`endif 

`ifdef i_axi_AXI_W_MCA_NC_W_S15
  `define AXI_W_MCA_NC_W_S15 `i_axi_AXI_W_MCA_NC_W_S15
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_S16
  `define AXI_AR_MCA_NC_S16 `i_axi_AXI_AR_MCA_NC_S16
`endif 

`ifdef i_axi_AXI_AR_MCA_EN_S16
  `define AXI_AR_MCA_EN_S16 `i_axi_AXI_AR_MCA_EN_S16
`endif 

`ifdef i_axi_AXI_AR_MCA_NC_W_S16
  `define AXI_AR_MCA_NC_W_S16 `i_axi_AXI_AR_MCA_NC_W_S16
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_S16
  `define AXI_AW_MCA_NC_S16 `i_axi_AXI_AW_MCA_NC_S16
`endif 

`ifdef i_axi_AXI_AW_MCA_EN_S16
  `define AXI_AW_MCA_EN_S16 `i_axi_AXI_AW_MCA_EN_S16
`endif 

`ifdef i_axi_AXI_AW_MCA_NC_W_S16
  `define AXI_AW_MCA_NC_W_S16 `i_axi_AXI_AW_MCA_NC_W_S16
`endif 

`ifdef i_axi_AXI_W_MCA_NC_S16
  `define AXI_W_MCA_NC_S16 `i_axi_AXI_W_MCA_NC_S16
`endif 

`ifdef i_axi_AXI_W_MCA_EN_S16
  `define AXI_W_MCA_EN_S16 `i_axi_AXI_W_MCA_EN_S16
`endif 

`ifdef i_axi_AXI_W_MCA_NC_W_S16
  `define AXI_W_MCA_NC_W_S16 `i_axi_AXI_W_MCA_NC_W_S16
`endif 

`ifdef i_axi_AXI_R_MCA_NC_M1
  `define AXI_R_MCA_NC_M1 `i_axi_AXI_R_MCA_NC_M1
`endif 

`ifdef i_axi_AXI_R_MCA_EN_M1
  `define AXI_R_MCA_EN_M1 `i_axi_AXI_R_MCA_EN_M1
`endif 

`ifdef i_axi_AXI_R_MCA_NC_W_M1
  `define AXI_R_MCA_NC_W_M1 `i_axi_AXI_R_MCA_NC_W_M1
`endif 

`ifdef i_axi_AXI_B_MCA_NC_M1
  `define AXI_B_MCA_NC_M1 `i_axi_AXI_B_MCA_NC_M1
`endif 

`ifdef i_axi_AXI_B_MCA_EN_M1
  `define AXI_B_MCA_EN_M1 `i_axi_AXI_B_MCA_EN_M1
`endif 

`ifdef i_axi_AXI_B_MCA_NC_W_M1
  `define AXI_B_MCA_NC_W_M1 `i_axi_AXI_B_MCA_NC_W_M1
`endif 

`ifdef i_axi_AXI_R_MCA_NC_M2
  `define AXI_R_MCA_NC_M2 `i_axi_AXI_R_MCA_NC_M2
`endif 

`ifdef i_axi_AXI_R_MCA_EN_M2
  `define AXI_R_MCA_EN_M2 `i_axi_AXI_R_MCA_EN_M2
`endif 

`ifdef i_axi_AXI_R_MCA_NC_W_M2
  `define AXI_R_MCA_NC_W_M2 `i_axi_AXI_R_MCA_NC_W_M2
`endif 

`ifdef i_axi_AXI_B_MCA_NC_M2
  `define AXI_B_MCA_NC_M2 `i_axi_AXI_B_MCA_NC_M2
`endif 

`ifdef i_axi_AXI_B_MCA_EN_M2
  `define AXI_B_MCA_EN_M2 `i_axi_AXI_B_MCA_EN_M2
`endif 

`ifdef i_axi_AXI_B_MCA_NC_W_M2
  `define AXI_B_MCA_NC_W_M2 `i_axi_AXI_B_MCA_NC_W_M2
`endif 

`ifdef i_axi_AXI_R_MCA_NC_M3
  `define AXI_R_MCA_NC_M3 `i_axi_AXI_R_MCA_NC_M3
`endif 

`ifdef i_axi_AXI_R_MCA_EN_M3
  `define AXI_R_MCA_EN_M3 `i_axi_AXI_R_MCA_EN_M3
`endif 

`ifdef i_axi_AXI_R_MCA_NC_W_M3
  `define AXI_R_MCA_NC_W_M3 `i_axi_AXI_R_MCA_NC_W_M3
`endif 

`ifdef i_axi_AXI_B_MCA_NC_M3
  `define AXI_B_MCA_NC_M3 `i_axi_AXI_B_MCA_NC_M3
`endif 

`ifdef i_axi_AXI_B_MCA_EN_M3
  `define AXI_B_MCA_EN_M3 `i_axi_AXI_B_MCA_EN_M3
`endif 

`ifdef i_axi_AXI_B_MCA_NC_W_M3
  `define AXI_B_MCA_NC_W_M3 `i_axi_AXI_B_MCA_NC_W_M3
`endif 

`ifdef i_axi_AXI_R_MCA_NC_M4
  `define AXI_R_MCA_NC_M4 `i_axi_AXI_R_MCA_NC_M4
`endif 

`ifdef i_axi_AXI_R_MCA_EN_M4
  `define AXI_R_MCA_EN_M4 `i_axi_AXI_R_MCA_EN_M4
`endif 

`ifdef i_axi_AXI_R_MCA_NC_W_M4
  `define AXI_R_MCA_NC_W_M4 `i_axi_AXI_R_MCA_NC_W_M4
`endif 

`ifdef i_axi_AXI_B_MCA_NC_M4
  `define AXI_B_MCA_NC_M4 `i_axi_AXI_B_MCA_NC_M4
`endif 

`ifdef i_axi_AXI_B_MCA_EN_M4
  `define AXI_B_MCA_EN_M4 `i_axi_AXI_B_MCA_EN_M4
`endif 

`ifdef i_axi_AXI_B_MCA_NC_W_M4
  `define AXI_B_MCA_NC_W_M4 `i_axi_AXI_B_MCA_NC_W_M4
`endif 

`ifdef i_axi_AXI_R_MCA_NC_M5
  `define AXI_R_MCA_NC_M5 `i_axi_AXI_R_MCA_NC_M5
`endif 

`ifdef i_axi_AXI_R_MCA_EN_M5
  `define AXI_R_MCA_EN_M5 `i_axi_AXI_R_MCA_EN_M5
`endif 

`ifdef i_axi_AXI_R_MCA_NC_W_M5
  `define AXI_R_MCA_NC_W_M5 `i_axi_AXI_R_MCA_NC_W_M5
`endif 

`ifdef i_axi_AXI_B_MCA_NC_M5
  `define AXI_B_MCA_NC_M5 `i_axi_AXI_B_MCA_NC_M5
`endif 

`ifdef i_axi_AXI_B_MCA_EN_M5
  `define AXI_B_MCA_EN_M5 `i_axi_AXI_B_MCA_EN_M5
`endif 

`ifdef i_axi_AXI_B_MCA_NC_W_M5
  `define AXI_B_MCA_NC_W_M5 `i_axi_AXI_B_MCA_NC_W_M5
`endif 

`ifdef i_axi_AXI_R_MCA_NC_M6
  `define AXI_R_MCA_NC_M6 `i_axi_AXI_R_MCA_NC_M6
`endif 

`ifdef i_axi_AXI_R_MCA_EN_M6
  `define AXI_R_MCA_EN_M6 `i_axi_AXI_R_MCA_EN_M6
`endif 

`ifdef i_axi_AXI_R_MCA_NC_W_M6
  `define AXI_R_MCA_NC_W_M6 `i_axi_AXI_R_MCA_NC_W_M6
`endif 

`ifdef i_axi_AXI_B_MCA_NC_M6
  `define AXI_B_MCA_NC_M6 `i_axi_AXI_B_MCA_NC_M6
`endif 

`ifdef i_axi_AXI_B_MCA_EN_M6
  `define AXI_B_MCA_EN_M6 `i_axi_AXI_B_MCA_EN_M6
`endif 

`ifdef i_axi_AXI_B_MCA_NC_W_M6
  `define AXI_B_MCA_NC_W_M6 `i_axi_AXI_B_MCA_NC_W_M6
`endif 

`ifdef i_axi_AXI_R_MCA_NC_M7
  `define AXI_R_MCA_NC_M7 `i_axi_AXI_R_MCA_NC_M7
`endif 

`ifdef i_axi_AXI_R_MCA_EN_M7
  `define AXI_R_MCA_EN_M7 `i_axi_AXI_R_MCA_EN_M7
`endif 

`ifdef i_axi_AXI_R_MCA_NC_W_M7
  `define AXI_R_MCA_NC_W_M7 `i_axi_AXI_R_MCA_NC_W_M7
`endif 

`ifdef i_axi_AXI_B_MCA_NC_M7
  `define AXI_B_MCA_NC_M7 `i_axi_AXI_B_MCA_NC_M7
`endif 

`ifdef i_axi_AXI_B_MCA_EN_M7
  `define AXI_B_MCA_EN_M7 `i_axi_AXI_B_MCA_EN_M7
`endif 

`ifdef i_axi_AXI_B_MCA_NC_W_M7
  `define AXI_B_MCA_NC_W_M7 `i_axi_AXI_B_MCA_NC_W_M7
`endif 

`ifdef i_axi_AXI_R_MCA_NC_M8
  `define AXI_R_MCA_NC_M8 `i_axi_AXI_R_MCA_NC_M8
`endif 

`ifdef i_axi_AXI_R_MCA_EN_M8
  `define AXI_R_MCA_EN_M8 `i_axi_AXI_R_MCA_EN_M8
`endif 

`ifdef i_axi_AXI_R_MCA_NC_W_M8
  `define AXI_R_MCA_NC_W_M8 `i_axi_AXI_R_MCA_NC_W_M8
`endif 

`ifdef i_axi_AXI_B_MCA_NC_M8
  `define AXI_B_MCA_NC_M8 `i_axi_AXI_B_MCA_NC_M8
`endif 

`ifdef i_axi_AXI_B_MCA_EN_M8
  `define AXI_B_MCA_EN_M8 `i_axi_AXI_B_MCA_EN_M8
`endif 

`ifdef i_axi_AXI_B_MCA_NC_W_M8
  `define AXI_B_MCA_NC_W_M8 `i_axi_AXI_B_MCA_NC_W_M8
`endif 

`ifdef i_axi_AXI_R_MCA_NC_M9
  `define AXI_R_MCA_NC_M9 `i_axi_AXI_R_MCA_NC_M9
`endif 

`ifdef i_axi_AXI_R_MCA_EN_M9
  `define AXI_R_MCA_EN_M9 `i_axi_AXI_R_MCA_EN_M9
`endif 

`ifdef i_axi_AXI_R_MCA_NC_W_M9
  `define AXI_R_MCA_NC_W_M9 `i_axi_AXI_R_MCA_NC_W_M9
`endif 

`ifdef i_axi_AXI_B_MCA_NC_M9
  `define AXI_B_MCA_NC_M9 `i_axi_AXI_B_MCA_NC_M9
`endif 

`ifdef i_axi_AXI_B_MCA_EN_M9
  `define AXI_B_MCA_EN_M9 `i_axi_AXI_B_MCA_EN_M9
`endif 

`ifdef i_axi_AXI_B_MCA_NC_W_M9
  `define AXI_B_MCA_NC_W_M9 `i_axi_AXI_B_MCA_NC_W_M9
`endif 

`ifdef i_axi_AXI_R_MCA_NC_M10
  `define AXI_R_MCA_NC_M10 `i_axi_AXI_R_MCA_NC_M10
`endif 

`ifdef i_axi_AXI_R_MCA_EN_M10
  `define AXI_R_MCA_EN_M10 `i_axi_AXI_R_MCA_EN_M10
`endif 

`ifdef i_axi_AXI_R_MCA_NC_W_M10
  `define AXI_R_MCA_NC_W_M10 `i_axi_AXI_R_MCA_NC_W_M10
`endif 

`ifdef i_axi_AXI_B_MCA_NC_M10
  `define AXI_B_MCA_NC_M10 `i_axi_AXI_B_MCA_NC_M10
`endif 

`ifdef i_axi_AXI_B_MCA_EN_M10
  `define AXI_B_MCA_EN_M10 `i_axi_AXI_B_MCA_EN_M10
`endif 

`ifdef i_axi_AXI_B_MCA_NC_W_M10
  `define AXI_B_MCA_NC_W_M10 `i_axi_AXI_B_MCA_NC_W_M10
`endif 

`ifdef i_axi_AXI_R_MCA_NC_M11
  `define AXI_R_MCA_NC_M11 `i_axi_AXI_R_MCA_NC_M11
`endif 

`ifdef i_axi_AXI_R_MCA_EN_M11
  `define AXI_R_MCA_EN_M11 `i_axi_AXI_R_MCA_EN_M11
`endif 

`ifdef i_axi_AXI_R_MCA_NC_W_M11
  `define AXI_R_MCA_NC_W_M11 `i_axi_AXI_R_MCA_NC_W_M11
`endif 

`ifdef i_axi_AXI_B_MCA_NC_M11
  `define AXI_B_MCA_NC_M11 `i_axi_AXI_B_MCA_NC_M11
`endif 

`ifdef i_axi_AXI_B_MCA_EN_M11
  `define AXI_B_MCA_EN_M11 `i_axi_AXI_B_MCA_EN_M11
`endif 

`ifdef i_axi_AXI_B_MCA_NC_W_M11
  `define AXI_B_MCA_NC_W_M11 `i_axi_AXI_B_MCA_NC_W_M11
`endif 

`ifdef i_axi_AXI_R_MCA_NC_M12
  `define AXI_R_MCA_NC_M12 `i_axi_AXI_R_MCA_NC_M12
`endif 

`ifdef i_axi_AXI_R_MCA_EN_M12
  `define AXI_R_MCA_EN_M12 `i_axi_AXI_R_MCA_EN_M12
`endif 

`ifdef i_axi_AXI_R_MCA_NC_W_M12
  `define AXI_R_MCA_NC_W_M12 `i_axi_AXI_R_MCA_NC_W_M12
`endif 

`ifdef i_axi_AXI_B_MCA_NC_M12
  `define AXI_B_MCA_NC_M12 `i_axi_AXI_B_MCA_NC_M12
`endif 

`ifdef i_axi_AXI_B_MCA_EN_M12
  `define AXI_B_MCA_EN_M12 `i_axi_AXI_B_MCA_EN_M12
`endif 

`ifdef i_axi_AXI_B_MCA_NC_W_M12
  `define AXI_B_MCA_NC_W_M12 `i_axi_AXI_B_MCA_NC_W_M12
`endif 

`ifdef i_axi_AXI_R_MCA_NC_M13
  `define AXI_R_MCA_NC_M13 `i_axi_AXI_R_MCA_NC_M13
`endif 

`ifdef i_axi_AXI_R_MCA_EN_M13
  `define AXI_R_MCA_EN_M13 `i_axi_AXI_R_MCA_EN_M13
`endif 

`ifdef i_axi_AXI_R_MCA_NC_W_M13
  `define AXI_R_MCA_NC_W_M13 `i_axi_AXI_R_MCA_NC_W_M13
`endif 

`ifdef i_axi_AXI_B_MCA_NC_M13
  `define AXI_B_MCA_NC_M13 `i_axi_AXI_B_MCA_NC_M13
`endif 

`ifdef i_axi_AXI_B_MCA_EN_M13
  `define AXI_B_MCA_EN_M13 `i_axi_AXI_B_MCA_EN_M13
`endif 

`ifdef i_axi_AXI_B_MCA_NC_W_M13
  `define AXI_B_MCA_NC_W_M13 `i_axi_AXI_B_MCA_NC_W_M13
`endif 

`ifdef i_axi_AXI_R_MCA_NC_M14
  `define AXI_R_MCA_NC_M14 `i_axi_AXI_R_MCA_NC_M14
`endif 

`ifdef i_axi_AXI_R_MCA_EN_M14
  `define AXI_R_MCA_EN_M14 `i_axi_AXI_R_MCA_EN_M14
`endif 

`ifdef i_axi_AXI_R_MCA_NC_W_M14
  `define AXI_R_MCA_NC_W_M14 `i_axi_AXI_R_MCA_NC_W_M14
`endif 

`ifdef i_axi_AXI_B_MCA_NC_M14
  `define AXI_B_MCA_NC_M14 `i_axi_AXI_B_MCA_NC_M14
`endif 

`ifdef i_axi_AXI_B_MCA_EN_M14
  `define AXI_B_MCA_EN_M14 `i_axi_AXI_B_MCA_EN_M14
`endif 

`ifdef i_axi_AXI_B_MCA_NC_W_M14
  `define AXI_B_MCA_NC_W_M14 `i_axi_AXI_B_MCA_NC_W_M14
`endif 

`ifdef i_axi_AXI_R_MCA_NC_M15
  `define AXI_R_MCA_NC_M15 `i_axi_AXI_R_MCA_NC_M15
`endif 

`ifdef i_axi_AXI_R_MCA_EN_M15
  `define AXI_R_MCA_EN_M15 `i_axi_AXI_R_MCA_EN_M15
`endif 

`ifdef i_axi_AXI_R_MCA_NC_W_M15
  `define AXI_R_MCA_NC_W_M15 `i_axi_AXI_R_MCA_NC_W_M15
`endif 

`ifdef i_axi_AXI_B_MCA_NC_M15
  `define AXI_B_MCA_NC_M15 `i_axi_AXI_B_MCA_NC_M15
`endif 

`ifdef i_axi_AXI_B_MCA_EN_M15
  `define AXI_B_MCA_EN_M15 `i_axi_AXI_B_MCA_EN_M15
`endif 

`ifdef i_axi_AXI_B_MCA_NC_W_M15
  `define AXI_B_MCA_NC_W_M15 `i_axi_AXI_B_MCA_NC_W_M15
`endif 

`ifdef i_axi_AXI_R_MCA_NC_M16
  `define AXI_R_MCA_NC_M16 `i_axi_AXI_R_MCA_NC_M16
`endif 

`ifdef i_axi_AXI_R_MCA_EN_M16
  `define AXI_R_MCA_EN_M16 `i_axi_AXI_R_MCA_EN_M16
`endif 

`ifdef i_axi_AXI_R_MCA_NC_W_M16
  `define AXI_R_MCA_NC_W_M16 `i_axi_AXI_R_MCA_NC_W_M16
`endif 

`ifdef i_axi_AXI_B_MCA_NC_M16
  `define AXI_B_MCA_NC_M16 `i_axi_AXI_B_MCA_NC_M16
`endif 

`ifdef i_axi_AXI_B_MCA_EN_M16
  `define AXI_B_MCA_EN_M16 `i_axi_AXI_B_MCA_EN_M16
`endif 

`ifdef i_axi_AXI_B_MCA_NC_W_M16
  `define AXI_B_MCA_NC_W_M16 `i_axi_AXI_B_MCA_NC_W_M16
`endif 

`ifdef i_axi_AXI_AR_SHARED_MCA_NC
  `define AXI_AR_SHARED_MCA_NC `i_axi_AXI_AR_SHARED_MCA_NC
`endif 

`ifdef i_axi_AXI_AR_SHARED_MCA_EN
  `define AXI_AR_SHARED_MCA_EN `i_axi_AXI_AR_SHARED_MCA_EN
`endif 

`ifdef i_axi_AXI_AR_SHARED_MCA_NC_W
  `define AXI_AR_SHARED_MCA_NC_W `i_axi_AXI_AR_SHARED_MCA_NC_W
`endif 

`ifdef i_axi_AXI_AW_SHARED_MCA_NC
  `define AXI_AW_SHARED_MCA_NC `i_axi_AXI_AW_SHARED_MCA_NC
`endif 

`ifdef i_axi_AXI_AW_SHARED_MCA_EN
  `define AXI_AW_SHARED_MCA_EN `i_axi_AXI_AW_SHARED_MCA_EN
`endif 

`ifdef i_axi_AXI_AW_SHARED_MCA_NC_W
  `define AXI_AW_SHARED_MCA_NC_W `i_axi_AXI_AW_SHARED_MCA_NC_W
`endif 

`ifdef i_axi_AXI_W_SHARED_MCA_NC
  `define AXI_W_SHARED_MCA_NC `i_axi_AXI_W_SHARED_MCA_NC
`endif 

`ifdef i_axi_AXI_W_SHARED_MCA_EN
  `define AXI_W_SHARED_MCA_EN `i_axi_AXI_W_SHARED_MCA_EN
`endif 

`ifdef i_axi_AXI_W_SHARED_MCA_NC_W
  `define AXI_W_SHARED_MCA_NC_W `i_axi_AXI_W_SHARED_MCA_NC_W
`endif 

`ifdef i_axi_AXI_R_SHARED_MCA_NC
  `define AXI_R_SHARED_MCA_NC `i_axi_AXI_R_SHARED_MCA_NC
`endif 

`ifdef i_axi_AXI_R_SHARED_MCA_EN
  `define AXI_R_SHARED_MCA_EN `i_axi_AXI_R_SHARED_MCA_EN
`endif 

`ifdef i_axi_AXI_R_SHARED_MCA_NC_W
  `define AXI_R_SHARED_MCA_NC_W `i_axi_AXI_R_SHARED_MCA_NC_W
`endif 

`ifdef i_axi_AXI_B_SHARED_MCA_NC
  `define AXI_B_SHARED_MCA_NC `i_axi_AXI_B_SHARED_MCA_NC
`endif 

`ifdef i_axi_AXI_B_SHARED_MCA_EN
  `define AXI_B_SHARED_MCA_EN `i_axi_AXI_B_SHARED_MCA_EN
`endif 

`ifdef i_axi_AXI_B_SHARED_MCA_NC_W
  `define AXI_B_SHARED_MCA_NC_W `i_axi_AXI_B_SHARED_MCA_NC_W
`endif 

`ifdef i_axi_AXI_MAX_RCA_ID_M1
  `define AXI_MAX_RCA_ID_M1 `i_axi_AXI_MAX_RCA_ID_M1
`endif 

`ifdef i_axi_AXI_LOG2_MAX_RCA_ID_P1_M1
  `define AXI_LOG2_MAX_RCA_ID_P1_M1 `i_axi_AXI_LOG2_MAX_RCA_ID_P1_M1
`endif 

`ifdef i_axi_AXI_MAX_WCA_ID_M1
  `define AXI_MAX_WCA_ID_M1 `i_axi_AXI_MAX_WCA_ID_M1
`endif 

`ifdef i_axi_AXI_LOG2_MAX_WCA_ID_P1_M1
  `define AXI_LOG2_MAX_WCA_ID_P1_M1 `i_axi_AXI_LOG2_MAX_WCA_ID_P1_M1
`endif 

`ifdef i_axi_AXI_MAX_URIDA_M1
  `define AXI_MAX_URIDA_M1 `i_axi_AXI_MAX_URIDA_M1
`endif 

`ifdef i_axi_AXI_LOG2_MAX_URIDA_M1
  `define AXI_LOG2_MAX_URIDA_M1 `i_axi_AXI_LOG2_MAX_URIDA_M1
`endif 

`ifdef i_axi_AXI_MAX_UWIDA_M1
  `define AXI_MAX_UWIDA_M1 `i_axi_AXI_MAX_UWIDA_M1
`endif 

`ifdef i_axi_AXI_LOG2_MAX_UWIDA_M1
  `define AXI_LOG2_MAX_UWIDA_M1 `i_axi_AXI_LOG2_MAX_UWIDA_M1
`endif 

`ifdef i_axi_AXI_RI_LIMIT_M1
  `define AXI_RI_LIMIT_M1 `i_axi_AXI_RI_LIMIT_M1
`endif 

`ifdef i_axi_AXI_MAX_RCA_ID_M2
  `define AXI_MAX_RCA_ID_M2 `i_axi_AXI_MAX_RCA_ID_M2
`endif 

`ifdef i_axi_AXI_LOG2_MAX_RCA_ID_P1_M2
  `define AXI_LOG2_MAX_RCA_ID_P1_M2 `i_axi_AXI_LOG2_MAX_RCA_ID_P1_M2
`endif 

`ifdef i_axi_AXI_MAX_WCA_ID_M2
  `define AXI_MAX_WCA_ID_M2 `i_axi_AXI_MAX_WCA_ID_M2
`endif 

`ifdef i_axi_AXI_LOG2_MAX_WCA_ID_P1_M2
  `define AXI_LOG2_MAX_WCA_ID_P1_M2 `i_axi_AXI_LOG2_MAX_WCA_ID_P1_M2
`endif 

`ifdef i_axi_AXI_MAX_URIDA_M2
  `define AXI_MAX_URIDA_M2 `i_axi_AXI_MAX_URIDA_M2
`endif 

`ifdef i_axi_AXI_LOG2_MAX_URIDA_M2
  `define AXI_LOG2_MAX_URIDA_M2 `i_axi_AXI_LOG2_MAX_URIDA_M2
`endif 

`ifdef i_axi_AXI_MAX_UWIDA_M2
  `define AXI_MAX_UWIDA_M2 `i_axi_AXI_MAX_UWIDA_M2
`endif 

`ifdef i_axi_AXI_LOG2_MAX_UWIDA_M2
  `define AXI_LOG2_MAX_UWIDA_M2 `i_axi_AXI_LOG2_MAX_UWIDA_M2
`endif 

`ifdef i_axi_AXI_RI_LIMIT_M2
  `define AXI_RI_LIMIT_M2 `i_axi_AXI_RI_LIMIT_M2
`endif 

`ifdef i_axi_AXI_MAX_RCA_ID_M3
  `define AXI_MAX_RCA_ID_M3 `i_axi_AXI_MAX_RCA_ID_M3
`endif 

`ifdef i_axi_AXI_LOG2_MAX_RCA_ID_P1_M3
  `define AXI_LOG2_MAX_RCA_ID_P1_M3 `i_axi_AXI_LOG2_MAX_RCA_ID_P1_M3
`endif 

`ifdef i_axi_AXI_MAX_WCA_ID_M3
  `define AXI_MAX_WCA_ID_M3 `i_axi_AXI_MAX_WCA_ID_M3
`endif 

`ifdef i_axi_AXI_LOG2_MAX_WCA_ID_P1_M3
  `define AXI_LOG2_MAX_WCA_ID_P1_M3 `i_axi_AXI_LOG2_MAX_WCA_ID_P1_M3
`endif 

`ifdef i_axi_AXI_MAX_URIDA_M3
  `define AXI_MAX_URIDA_M3 `i_axi_AXI_MAX_URIDA_M3
`endif 

`ifdef i_axi_AXI_LOG2_MAX_URIDA_M3
  `define AXI_LOG2_MAX_URIDA_M3 `i_axi_AXI_LOG2_MAX_URIDA_M3
`endif 

`ifdef i_axi_AXI_MAX_UWIDA_M3
  `define AXI_MAX_UWIDA_M3 `i_axi_AXI_MAX_UWIDA_M3
`endif 

`ifdef i_axi_AXI_LOG2_MAX_UWIDA_M3
  `define AXI_LOG2_MAX_UWIDA_M3 `i_axi_AXI_LOG2_MAX_UWIDA_M3
`endif 

`ifdef i_axi_AXI_RI_LIMIT_M3
  `define AXI_RI_LIMIT_M3 `i_axi_AXI_RI_LIMIT_M3
`endif 

`ifdef i_axi_AXI_MAX_RCA_ID_M4
  `define AXI_MAX_RCA_ID_M4 `i_axi_AXI_MAX_RCA_ID_M4
`endif 

`ifdef i_axi_AXI_LOG2_MAX_RCA_ID_P1_M4
  `define AXI_LOG2_MAX_RCA_ID_P1_M4 `i_axi_AXI_LOG2_MAX_RCA_ID_P1_M4
`endif 

`ifdef i_axi_AXI_MAX_WCA_ID_M4
  `define AXI_MAX_WCA_ID_M4 `i_axi_AXI_MAX_WCA_ID_M4
`endif 

`ifdef i_axi_AXI_LOG2_MAX_WCA_ID_P1_M4
  `define AXI_LOG2_MAX_WCA_ID_P1_M4 `i_axi_AXI_LOG2_MAX_WCA_ID_P1_M4
`endif 

`ifdef i_axi_AXI_MAX_URIDA_M4
  `define AXI_MAX_URIDA_M4 `i_axi_AXI_MAX_URIDA_M4
`endif 

`ifdef i_axi_AXI_LOG2_MAX_URIDA_M4
  `define AXI_LOG2_MAX_URIDA_M4 `i_axi_AXI_LOG2_MAX_URIDA_M4
`endif 

`ifdef i_axi_AXI_MAX_UWIDA_M4
  `define AXI_MAX_UWIDA_M4 `i_axi_AXI_MAX_UWIDA_M4
`endif 

`ifdef i_axi_AXI_LOG2_MAX_UWIDA_M4
  `define AXI_LOG2_MAX_UWIDA_M4 `i_axi_AXI_LOG2_MAX_UWIDA_M4
`endif 

`ifdef i_axi_AXI_RI_LIMIT_M4
  `define AXI_RI_LIMIT_M4 `i_axi_AXI_RI_LIMIT_M4
`endif 

`ifdef i_axi_AXI_MAX_RCA_ID_M5
  `define AXI_MAX_RCA_ID_M5 `i_axi_AXI_MAX_RCA_ID_M5
`endif 

`ifdef i_axi_AXI_LOG2_MAX_RCA_ID_P1_M5
  `define AXI_LOG2_MAX_RCA_ID_P1_M5 `i_axi_AXI_LOG2_MAX_RCA_ID_P1_M5
`endif 

`ifdef i_axi_AXI_MAX_WCA_ID_M5
  `define AXI_MAX_WCA_ID_M5 `i_axi_AXI_MAX_WCA_ID_M5
`endif 

`ifdef i_axi_AXI_LOG2_MAX_WCA_ID_P1_M5
  `define AXI_LOG2_MAX_WCA_ID_P1_M5 `i_axi_AXI_LOG2_MAX_WCA_ID_P1_M5
`endif 

`ifdef i_axi_AXI_MAX_URIDA_M5
  `define AXI_MAX_URIDA_M5 `i_axi_AXI_MAX_URIDA_M5
`endif 

`ifdef i_axi_AXI_LOG2_MAX_URIDA_M5
  `define AXI_LOG2_MAX_URIDA_M5 `i_axi_AXI_LOG2_MAX_URIDA_M5
`endif 

`ifdef i_axi_AXI_MAX_UWIDA_M5
  `define AXI_MAX_UWIDA_M5 `i_axi_AXI_MAX_UWIDA_M5
`endif 

`ifdef i_axi_AXI_LOG2_MAX_UWIDA_M5
  `define AXI_LOG2_MAX_UWIDA_M5 `i_axi_AXI_LOG2_MAX_UWIDA_M5
`endif 

`ifdef i_axi_AXI_RI_LIMIT_M5
  `define AXI_RI_LIMIT_M5 `i_axi_AXI_RI_LIMIT_M5
`endif 

`ifdef i_axi_AXI_MAX_RCA_ID_M6
  `define AXI_MAX_RCA_ID_M6 `i_axi_AXI_MAX_RCA_ID_M6
`endif 

`ifdef i_axi_AXI_LOG2_MAX_RCA_ID_P1_M6
  `define AXI_LOG2_MAX_RCA_ID_P1_M6 `i_axi_AXI_LOG2_MAX_RCA_ID_P1_M6
`endif 

`ifdef i_axi_AXI_MAX_WCA_ID_M6
  `define AXI_MAX_WCA_ID_M6 `i_axi_AXI_MAX_WCA_ID_M6
`endif 

`ifdef i_axi_AXI_LOG2_MAX_WCA_ID_P1_M6
  `define AXI_LOG2_MAX_WCA_ID_P1_M6 `i_axi_AXI_LOG2_MAX_WCA_ID_P1_M6
`endif 

`ifdef i_axi_AXI_MAX_URIDA_M6
  `define AXI_MAX_URIDA_M6 `i_axi_AXI_MAX_URIDA_M6
`endif 

`ifdef i_axi_AXI_LOG2_MAX_URIDA_M6
  `define AXI_LOG2_MAX_URIDA_M6 `i_axi_AXI_LOG2_MAX_URIDA_M6
`endif 

`ifdef i_axi_AXI_MAX_UWIDA_M6
  `define AXI_MAX_UWIDA_M6 `i_axi_AXI_MAX_UWIDA_M6
`endif 

`ifdef i_axi_AXI_LOG2_MAX_UWIDA_M6
  `define AXI_LOG2_MAX_UWIDA_M6 `i_axi_AXI_LOG2_MAX_UWIDA_M6
`endif 

`ifdef i_axi_AXI_RI_LIMIT_M6
  `define AXI_RI_LIMIT_M6 `i_axi_AXI_RI_LIMIT_M6
`endif 

`ifdef i_axi_AXI_MAX_RCA_ID_M7
  `define AXI_MAX_RCA_ID_M7 `i_axi_AXI_MAX_RCA_ID_M7
`endif 

`ifdef i_axi_AXI_LOG2_MAX_RCA_ID_P1_M7
  `define AXI_LOG2_MAX_RCA_ID_P1_M7 `i_axi_AXI_LOG2_MAX_RCA_ID_P1_M7
`endif 

`ifdef i_axi_AXI_MAX_WCA_ID_M7
  `define AXI_MAX_WCA_ID_M7 `i_axi_AXI_MAX_WCA_ID_M7
`endif 

`ifdef i_axi_AXI_LOG2_MAX_WCA_ID_P1_M7
  `define AXI_LOG2_MAX_WCA_ID_P1_M7 `i_axi_AXI_LOG2_MAX_WCA_ID_P1_M7
`endif 

`ifdef i_axi_AXI_MAX_URIDA_M7
  `define AXI_MAX_URIDA_M7 `i_axi_AXI_MAX_URIDA_M7
`endif 

`ifdef i_axi_AXI_LOG2_MAX_URIDA_M7
  `define AXI_LOG2_MAX_URIDA_M7 `i_axi_AXI_LOG2_MAX_URIDA_M7
`endif 

`ifdef i_axi_AXI_MAX_UWIDA_M7
  `define AXI_MAX_UWIDA_M7 `i_axi_AXI_MAX_UWIDA_M7
`endif 

`ifdef i_axi_AXI_LOG2_MAX_UWIDA_M7
  `define AXI_LOG2_MAX_UWIDA_M7 `i_axi_AXI_LOG2_MAX_UWIDA_M7
`endif 

`ifdef i_axi_AXI_RI_LIMIT_M7
  `define AXI_RI_LIMIT_M7 `i_axi_AXI_RI_LIMIT_M7
`endif 

`ifdef i_axi_AXI_MAX_RCA_ID_M8
  `define AXI_MAX_RCA_ID_M8 `i_axi_AXI_MAX_RCA_ID_M8
`endif 

`ifdef i_axi_AXI_LOG2_MAX_RCA_ID_P1_M8
  `define AXI_LOG2_MAX_RCA_ID_P1_M8 `i_axi_AXI_LOG2_MAX_RCA_ID_P1_M8
`endif 

`ifdef i_axi_AXI_MAX_WCA_ID_M8
  `define AXI_MAX_WCA_ID_M8 `i_axi_AXI_MAX_WCA_ID_M8
`endif 

`ifdef i_axi_AXI_LOG2_MAX_WCA_ID_P1_M8
  `define AXI_LOG2_MAX_WCA_ID_P1_M8 `i_axi_AXI_LOG2_MAX_WCA_ID_P1_M8
`endif 

`ifdef i_axi_AXI_MAX_URIDA_M8
  `define AXI_MAX_URIDA_M8 `i_axi_AXI_MAX_URIDA_M8
`endif 

`ifdef i_axi_AXI_LOG2_MAX_URIDA_M8
  `define AXI_LOG2_MAX_URIDA_M8 `i_axi_AXI_LOG2_MAX_URIDA_M8
`endif 

`ifdef i_axi_AXI_MAX_UWIDA_M8
  `define AXI_MAX_UWIDA_M8 `i_axi_AXI_MAX_UWIDA_M8
`endif 

`ifdef i_axi_AXI_LOG2_MAX_UWIDA_M8
  `define AXI_LOG2_MAX_UWIDA_M8 `i_axi_AXI_LOG2_MAX_UWIDA_M8
`endif 

`ifdef i_axi_AXI_RI_LIMIT_M8
  `define AXI_RI_LIMIT_M8 `i_axi_AXI_RI_LIMIT_M8
`endif 

`ifdef i_axi_AXI_MAX_RCA_ID_M9
  `define AXI_MAX_RCA_ID_M9 `i_axi_AXI_MAX_RCA_ID_M9
`endif 

`ifdef i_axi_AXI_LOG2_MAX_RCA_ID_P1_M9
  `define AXI_LOG2_MAX_RCA_ID_P1_M9 `i_axi_AXI_LOG2_MAX_RCA_ID_P1_M9
`endif 

`ifdef i_axi_AXI_MAX_WCA_ID_M9
  `define AXI_MAX_WCA_ID_M9 `i_axi_AXI_MAX_WCA_ID_M9
`endif 

`ifdef i_axi_AXI_LOG2_MAX_WCA_ID_P1_M9
  `define AXI_LOG2_MAX_WCA_ID_P1_M9 `i_axi_AXI_LOG2_MAX_WCA_ID_P1_M9
`endif 

`ifdef i_axi_AXI_MAX_URIDA_M9
  `define AXI_MAX_URIDA_M9 `i_axi_AXI_MAX_URIDA_M9
`endif 

`ifdef i_axi_AXI_LOG2_MAX_URIDA_M9
  `define AXI_LOG2_MAX_URIDA_M9 `i_axi_AXI_LOG2_MAX_URIDA_M9
`endif 

`ifdef i_axi_AXI_MAX_UWIDA_M9
  `define AXI_MAX_UWIDA_M9 `i_axi_AXI_MAX_UWIDA_M9
`endif 

`ifdef i_axi_AXI_LOG2_MAX_UWIDA_M9
  `define AXI_LOG2_MAX_UWIDA_M9 `i_axi_AXI_LOG2_MAX_UWIDA_M9
`endif 

`ifdef i_axi_AXI_RI_LIMIT_M9
  `define AXI_RI_LIMIT_M9 `i_axi_AXI_RI_LIMIT_M9
`endif 

`ifdef i_axi_AXI_MAX_RCA_ID_M10
  `define AXI_MAX_RCA_ID_M10 `i_axi_AXI_MAX_RCA_ID_M10
`endif 

`ifdef i_axi_AXI_LOG2_MAX_RCA_ID_P1_M10
  `define AXI_LOG2_MAX_RCA_ID_P1_M10 `i_axi_AXI_LOG2_MAX_RCA_ID_P1_M10
`endif 

`ifdef i_axi_AXI_MAX_WCA_ID_M10
  `define AXI_MAX_WCA_ID_M10 `i_axi_AXI_MAX_WCA_ID_M10
`endif 

`ifdef i_axi_AXI_LOG2_MAX_WCA_ID_P1_M10
  `define AXI_LOG2_MAX_WCA_ID_P1_M10 `i_axi_AXI_LOG2_MAX_WCA_ID_P1_M10
`endif 

`ifdef i_axi_AXI_MAX_URIDA_M10
  `define AXI_MAX_URIDA_M10 `i_axi_AXI_MAX_URIDA_M10
`endif 

`ifdef i_axi_AXI_LOG2_MAX_URIDA_M10
  `define AXI_LOG2_MAX_URIDA_M10 `i_axi_AXI_LOG2_MAX_URIDA_M10
`endif 

`ifdef i_axi_AXI_MAX_UWIDA_M10
  `define AXI_MAX_UWIDA_M10 `i_axi_AXI_MAX_UWIDA_M10
`endif 

`ifdef i_axi_AXI_LOG2_MAX_UWIDA_M10
  `define AXI_LOG2_MAX_UWIDA_M10 `i_axi_AXI_LOG2_MAX_UWIDA_M10
`endif 

`ifdef i_axi_AXI_RI_LIMIT_M10
  `define AXI_RI_LIMIT_M10 `i_axi_AXI_RI_LIMIT_M10
`endif 

`ifdef i_axi_AXI_MAX_RCA_ID_M11
  `define AXI_MAX_RCA_ID_M11 `i_axi_AXI_MAX_RCA_ID_M11
`endif 

`ifdef i_axi_AXI_LOG2_MAX_RCA_ID_P1_M11
  `define AXI_LOG2_MAX_RCA_ID_P1_M11 `i_axi_AXI_LOG2_MAX_RCA_ID_P1_M11
`endif 

`ifdef i_axi_AXI_MAX_WCA_ID_M11
  `define AXI_MAX_WCA_ID_M11 `i_axi_AXI_MAX_WCA_ID_M11
`endif 

`ifdef i_axi_AXI_LOG2_MAX_WCA_ID_P1_M11
  `define AXI_LOG2_MAX_WCA_ID_P1_M11 `i_axi_AXI_LOG2_MAX_WCA_ID_P1_M11
`endif 

`ifdef i_axi_AXI_MAX_URIDA_M11
  `define AXI_MAX_URIDA_M11 `i_axi_AXI_MAX_URIDA_M11
`endif 

`ifdef i_axi_AXI_LOG2_MAX_URIDA_M11
  `define AXI_LOG2_MAX_URIDA_M11 `i_axi_AXI_LOG2_MAX_URIDA_M11
`endif 

`ifdef i_axi_AXI_MAX_UWIDA_M11
  `define AXI_MAX_UWIDA_M11 `i_axi_AXI_MAX_UWIDA_M11
`endif 

`ifdef i_axi_AXI_LOG2_MAX_UWIDA_M11
  `define AXI_LOG2_MAX_UWIDA_M11 `i_axi_AXI_LOG2_MAX_UWIDA_M11
`endif 

`ifdef i_axi_AXI_RI_LIMIT_M11
  `define AXI_RI_LIMIT_M11 `i_axi_AXI_RI_LIMIT_M11
`endif 

`ifdef i_axi_AXI_MAX_RCA_ID_M12
  `define AXI_MAX_RCA_ID_M12 `i_axi_AXI_MAX_RCA_ID_M12
`endif 

`ifdef i_axi_AXI_LOG2_MAX_RCA_ID_P1_M12
  `define AXI_LOG2_MAX_RCA_ID_P1_M12 `i_axi_AXI_LOG2_MAX_RCA_ID_P1_M12
`endif 

`ifdef i_axi_AXI_MAX_WCA_ID_M12
  `define AXI_MAX_WCA_ID_M12 `i_axi_AXI_MAX_WCA_ID_M12
`endif 

`ifdef i_axi_AXI_LOG2_MAX_WCA_ID_P1_M12
  `define AXI_LOG2_MAX_WCA_ID_P1_M12 `i_axi_AXI_LOG2_MAX_WCA_ID_P1_M12
`endif 

`ifdef i_axi_AXI_MAX_URIDA_M12
  `define AXI_MAX_URIDA_M12 `i_axi_AXI_MAX_URIDA_M12
`endif 

`ifdef i_axi_AXI_LOG2_MAX_URIDA_M12
  `define AXI_LOG2_MAX_URIDA_M12 `i_axi_AXI_LOG2_MAX_URIDA_M12
`endif 

`ifdef i_axi_AXI_MAX_UWIDA_M12
  `define AXI_MAX_UWIDA_M12 `i_axi_AXI_MAX_UWIDA_M12
`endif 

`ifdef i_axi_AXI_LOG2_MAX_UWIDA_M12
  `define AXI_LOG2_MAX_UWIDA_M12 `i_axi_AXI_LOG2_MAX_UWIDA_M12
`endif 

`ifdef i_axi_AXI_RI_LIMIT_M12
  `define AXI_RI_LIMIT_M12 `i_axi_AXI_RI_LIMIT_M12
`endif 

`ifdef i_axi_AXI_MAX_RCA_ID_M13
  `define AXI_MAX_RCA_ID_M13 `i_axi_AXI_MAX_RCA_ID_M13
`endif 

`ifdef i_axi_AXI_LOG2_MAX_RCA_ID_P1_M13
  `define AXI_LOG2_MAX_RCA_ID_P1_M13 `i_axi_AXI_LOG2_MAX_RCA_ID_P1_M13
`endif 

`ifdef i_axi_AXI_MAX_WCA_ID_M13
  `define AXI_MAX_WCA_ID_M13 `i_axi_AXI_MAX_WCA_ID_M13
`endif 

`ifdef i_axi_AXI_LOG2_MAX_WCA_ID_P1_M13
  `define AXI_LOG2_MAX_WCA_ID_P1_M13 `i_axi_AXI_LOG2_MAX_WCA_ID_P1_M13
`endif 

`ifdef i_axi_AXI_MAX_URIDA_M13
  `define AXI_MAX_URIDA_M13 `i_axi_AXI_MAX_URIDA_M13
`endif 

`ifdef i_axi_AXI_LOG2_MAX_URIDA_M13
  `define AXI_LOG2_MAX_URIDA_M13 `i_axi_AXI_LOG2_MAX_URIDA_M13
`endif 

`ifdef i_axi_AXI_MAX_UWIDA_M13
  `define AXI_MAX_UWIDA_M13 `i_axi_AXI_MAX_UWIDA_M13
`endif 

`ifdef i_axi_AXI_LOG2_MAX_UWIDA_M13
  `define AXI_LOG2_MAX_UWIDA_M13 `i_axi_AXI_LOG2_MAX_UWIDA_M13
`endif 

`ifdef i_axi_AXI_RI_LIMIT_M13
  `define AXI_RI_LIMIT_M13 `i_axi_AXI_RI_LIMIT_M13
`endif 

`ifdef i_axi_AXI_MAX_RCA_ID_M14
  `define AXI_MAX_RCA_ID_M14 `i_axi_AXI_MAX_RCA_ID_M14
`endif 

`ifdef i_axi_AXI_LOG2_MAX_RCA_ID_P1_M14
  `define AXI_LOG2_MAX_RCA_ID_P1_M14 `i_axi_AXI_LOG2_MAX_RCA_ID_P1_M14
`endif 

`ifdef i_axi_AXI_MAX_WCA_ID_M14
  `define AXI_MAX_WCA_ID_M14 `i_axi_AXI_MAX_WCA_ID_M14
`endif 

`ifdef i_axi_AXI_LOG2_MAX_WCA_ID_P1_M14
  `define AXI_LOG2_MAX_WCA_ID_P1_M14 `i_axi_AXI_LOG2_MAX_WCA_ID_P1_M14
`endif 

`ifdef i_axi_AXI_MAX_URIDA_M14
  `define AXI_MAX_URIDA_M14 `i_axi_AXI_MAX_URIDA_M14
`endif 

`ifdef i_axi_AXI_LOG2_MAX_URIDA_M14
  `define AXI_LOG2_MAX_URIDA_M14 `i_axi_AXI_LOG2_MAX_URIDA_M14
`endif 

`ifdef i_axi_AXI_MAX_UWIDA_M14
  `define AXI_MAX_UWIDA_M14 `i_axi_AXI_MAX_UWIDA_M14
`endif 

`ifdef i_axi_AXI_LOG2_MAX_UWIDA_M14
  `define AXI_LOG2_MAX_UWIDA_M14 `i_axi_AXI_LOG2_MAX_UWIDA_M14
`endif 

`ifdef i_axi_AXI_RI_LIMIT_M14
  `define AXI_RI_LIMIT_M14 `i_axi_AXI_RI_LIMIT_M14
`endif 

`ifdef i_axi_AXI_MAX_RCA_ID_M15
  `define AXI_MAX_RCA_ID_M15 `i_axi_AXI_MAX_RCA_ID_M15
`endif 

`ifdef i_axi_AXI_LOG2_MAX_RCA_ID_P1_M15
  `define AXI_LOG2_MAX_RCA_ID_P1_M15 `i_axi_AXI_LOG2_MAX_RCA_ID_P1_M15
`endif 

`ifdef i_axi_AXI_MAX_WCA_ID_M15
  `define AXI_MAX_WCA_ID_M15 `i_axi_AXI_MAX_WCA_ID_M15
`endif 

`ifdef i_axi_AXI_LOG2_MAX_WCA_ID_P1_M15
  `define AXI_LOG2_MAX_WCA_ID_P1_M15 `i_axi_AXI_LOG2_MAX_WCA_ID_P1_M15
`endif 

`ifdef i_axi_AXI_MAX_URIDA_M15
  `define AXI_MAX_URIDA_M15 `i_axi_AXI_MAX_URIDA_M15
`endif 

`ifdef i_axi_AXI_LOG2_MAX_URIDA_M15
  `define AXI_LOG2_MAX_URIDA_M15 `i_axi_AXI_LOG2_MAX_URIDA_M15
`endif 

`ifdef i_axi_AXI_MAX_UWIDA_M15
  `define AXI_MAX_UWIDA_M15 `i_axi_AXI_MAX_UWIDA_M15
`endif 

`ifdef i_axi_AXI_LOG2_MAX_UWIDA_M15
  `define AXI_LOG2_MAX_UWIDA_M15 `i_axi_AXI_LOG2_MAX_UWIDA_M15
`endif 

`ifdef i_axi_AXI_RI_LIMIT_M15
  `define AXI_RI_LIMIT_M15 `i_axi_AXI_RI_LIMIT_M15
`endif 

`ifdef i_axi_AXI_MAX_RCA_ID_M16
  `define AXI_MAX_RCA_ID_M16 `i_axi_AXI_MAX_RCA_ID_M16
`endif 

`ifdef i_axi_AXI_LOG2_MAX_RCA_ID_P1_M16
  `define AXI_LOG2_MAX_RCA_ID_P1_M16 `i_axi_AXI_LOG2_MAX_RCA_ID_P1_M16
`endif 

`ifdef i_axi_AXI_MAX_WCA_ID_M16
  `define AXI_MAX_WCA_ID_M16 `i_axi_AXI_MAX_WCA_ID_M16
`endif 

`ifdef i_axi_AXI_LOG2_MAX_WCA_ID_P1_M16
  `define AXI_LOG2_MAX_WCA_ID_P1_M16 `i_axi_AXI_LOG2_MAX_WCA_ID_P1_M16
`endif 

`ifdef i_axi_AXI_MAX_URIDA_M16
  `define AXI_MAX_URIDA_M16 `i_axi_AXI_MAX_URIDA_M16
`endif 

`ifdef i_axi_AXI_LOG2_MAX_URIDA_M16
  `define AXI_LOG2_MAX_URIDA_M16 `i_axi_AXI_LOG2_MAX_URIDA_M16
`endif 

`ifdef i_axi_AXI_MAX_UWIDA_M16
  `define AXI_MAX_UWIDA_M16 `i_axi_AXI_MAX_UWIDA_M16
`endif 

`ifdef i_axi_AXI_LOG2_MAX_UWIDA_M16
  `define AXI_LOG2_MAX_UWIDA_M16 `i_axi_AXI_LOG2_MAX_UWIDA_M16
`endif 

`ifdef i_axi_AXI_RI_LIMIT_M16
  `define AXI_RI_LIMIT_M16 `i_axi_AXI_RI_LIMIT_M16
`endif 

`ifdef i_axi_AXI_MAX_FAWC_S0
  `define AXI_MAX_FAWC_S0 `i_axi_AXI_MAX_FAWC_S0
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_S0
  `define AXI_LOG2_MAX_FAWC_S0 `i_axi_AXI_LOG2_MAX_FAWC_S0
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_P1_S0
  `define AXI_LOG2_MAX_FAWC_P1_S0 `i_axi_AXI_LOG2_MAX_FAWC_P1_S0
`endif 

`ifdef i_axi_AXI_MAX_FARC_S0
  `define AXI_MAX_FARC_S0 `i_axi_AXI_MAX_FARC_S0
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FARC_P1_S0
  `define AXI_LOG2_MAX_FARC_P1_S0 `i_axi_AXI_LOG2_MAX_FARC_P1_S0
`endif 

`ifdef i_axi_AXI_WID_S0
  `define AXI_WID_S0 `i_axi_AXI_WID_S0
`endif 

`ifdef i_axi_AXI_MAX_FAC_EN
  `define AXI_MAX_FAC_EN `i_axi_AXI_MAX_FAC_EN
`endif 

`ifdef i_axi_AXI_WID_S1
  `define AXI_WID_S1 `i_axi_AXI_WID_S1
`endif 

`ifdef i_axi_AXI_LOG2_WID_S1
  `define AXI_LOG2_WID_S1 `i_axi_AXI_LOG2_WID_S1
`endif 

`ifdef i_axi_AXI_LOG2_WID_P1_S1
  `define AXI_LOG2_WID_P1_S1 `i_axi_AXI_LOG2_WID_P1_S1
`endif 

`ifdef i_axi_AXI_MAX_FAWC_S1
  `define AXI_MAX_FAWC_S1 `i_axi_AXI_MAX_FAWC_S1
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_S1
  `define AXI_LOG2_MAX_FAWC_S1 `i_axi_AXI_LOG2_MAX_FAWC_S1
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_P1_S1
  `define AXI_LOG2_MAX_FAWC_P1_S1 `i_axi_AXI_LOG2_MAX_FAWC_P1_S1
`endif 

`ifdef i_axi_AXI_MAX_FARC_S1
  `define AXI_MAX_FARC_S1 `i_axi_AXI_MAX_FARC_S1
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FARC_P1_S1
  `define AXI_LOG2_MAX_FARC_P1_S1 `i_axi_AXI_LOG2_MAX_FARC_P1_S1
`endif 

`ifdef i_axi_AXI_WID_S2
  `define AXI_WID_S2 `i_axi_AXI_WID_S2
`endif 

`ifdef i_axi_AXI_LOG2_WID_S2
  `define AXI_LOG2_WID_S2 `i_axi_AXI_LOG2_WID_S2
`endif 

`ifdef i_axi_AXI_LOG2_WID_P1_S2
  `define AXI_LOG2_WID_P1_S2 `i_axi_AXI_LOG2_WID_P1_S2
`endif 

`ifdef i_axi_AXI_MAX_FAWC_S2
  `define AXI_MAX_FAWC_S2 `i_axi_AXI_MAX_FAWC_S2
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_S2
  `define AXI_LOG2_MAX_FAWC_S2 `i_axi_AXI_LOG2_MAX_FAWC_S2
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_P1_S2
  `define AXI_LOG2_MAX_FAWC_P1_S2 `i_axi_AXI_LOG2_MAX_FAWC_P1_S2
`endif 

`ifdef i_axi_AXI_MAX_FARC_S2
  `define AXI_MAX_FARC_S2 `i_axi_AXI_MAX_FARC_S2
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FARC_P1_S2
  `define AXI_LOG2_MAX_FARC_P1_S2 `i_axi_AXI_LOG2_MAX_FARC_P1_S2
`endif 

`ifdef i_axi_AXI_WID_S3
  `define AXI_WID_S3 `i_axi_AXI_WID_S3
`endif 

`ifdef i_axi_AXI_LOG2_WID_S3
  `define AXI_LOG2_WID_S3 `i_axi_AXI_LOG2_WID_S3
`endif 

`ifdef i_axi_AXI_LOG2_WID_P1_S3
  `define AXI_LOG2_WID_P1_S3 `i_axi_AXI_LOG2_WID_P1_S3
`endif 

`ifdef i_axi_AXI_MAX_FAWC_S3
  `define AXI_MAX_FAWC_S3 `i_axi_AXI_MAX_FAWC_S3
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_S3
  `define AXI_LOG2_MAX_FAWC_S3 `i_axi_AXI_LOG2_MAX_FAWC_S3
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_P1_S3
  `define AXI_LOG2_MAX_FAWC_P1_S3 `i_axi_AXI_LOG2_MAX_FAWC_P1_S3
`endif 

`ifdef i_axi_AXI_MAX_FARC_S3
  `define AXI_MAX_FARC_S3 `i_axi_AXI_MAX_FARC_S3
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FARC_P1_S3
  `define AXI_LOG2_MAX_FARC_P1_S3 `i_axi_AXI_LOG2_MAX_FARC_P1_S3
`endif 

`ifdef i_axi_AXI_WID_S4
  `define AXI_WID_S4 `i_axi_AXI_WID_S4
`endif 

`ifdef i_axi_AXI_LOG2_WID_S4
  `define AXI_LOG2_WID_S4 `i_axi_AXI_LOG2_WID_S4
`endif 

`ifdef i_axi_AXI_LOG2_WID_P1_S4
  `define AXI_LOG2_WID_P1_S4 `i_axi_AXI_LOG2_WID_P1_S4
`endif 

`ifdef i_axi_AXI_MAX_FAWC_S4
  `define AXI_MAX_FAWC_S4 `i_axi_AXI_MAX_FAWC_S4
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_S4
  `define AXI_LOG2_MAX_FAWC_S4 `i_axi_AXI_LOG2_MAX_FAWC_S4
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_P1_S4
  `define AXI_LOG2_MAX_FAWC_P1_S4 `i_axi_AXI_LOG2_MAX_FAWC_P1_S4
`endif 

`ifdef i_axi_AXI_MAX_FARC_S4
  `define AXI_MAX_FARC_S4 `i_axi_AXI_MAX_FARC_S4
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FARC_P1_S4
  `define AXI_LOG2_MAX_FARC_P1_S4 `i_axi_AXI_LOG2_MAX_FARC_P1_S4
`endif 

`ifdef i_axi_AXI_WID_S5
  `define AXI_WID_S5 `i_axi_AXI_WID_S5
`endif 

`ifdef i_axi_AXI_LOG2_WID_S5
  `define AXI_LOG2_WID_S5 `i_axi_AXI_LOG2_WID_S5
`endif 

`ifdef i_axi_AXI_LOG2_WID_P1_S5
  `define AXI_LOG2_WID_P1_S5 `i_axi_AXI_LOG2_WID_P1_S5
`endif 

`ifdef i_axi_AXI_MAX_FAWC_S5
  `define AXI_MAX_FAWC_S5 `i_axi_AXI_MAX_FAWC_S5
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_S5
  `define AXI_LOG2_MAX_FAWC_S5 `i_axi_AXI_LOG2_MAX_FAWC_S5
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_P1_S5
  `define AXI_LOG2_MAX_FAWC_P1_S5 `i_axi_AXI_LOG2_MAX_FAWC_P1_S5
`endif 

`ifdef i_axi_AXI_MAX_FARC_S5
  `define AXI_MAX_FARC_S5 `i_axi_AXI_MAX_FARC_S5
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FARC_P1_S5
  `define AXI_LOG2_MAX_FARC_P1_S5 `i_axi_AXI_LOG2_MAX_FARC_P1_S5
`endif 

`ifdef i_axi_AXI_WID_S6
  `define AXI_WID_S6 `i_axi_AXI_WID_S6
`endif 

`ifdef i_axi_AXI_LOG2_WID_S6
  `define AXI_LOG2_WID_S6 `i_axi_AXI_LOG2_WID_S6
`endif 

`ifdef i_axi_AXI_LOG2_WID_P1_S6
  `define AXI_LOG2_WID_P1_S6 `i_axi_AXI_LOG2_WID_P1_S6
`endif 

`ifdef i_axi_AXI_MAX_FAWC_S6
  `define AXI_MAX_FAWC_S6 `i_axi_AXI_MAX_FAWC_S6
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_S6
  `define AXI_LOG2_MAX_FAWC_S6 `i_axi_AXI_LOG2_MAX_FAWC_S6
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_P1_S6
  `define AXI_LOG2_MAX_FAWC_P1_S6 `i_axi_AXI_LOG2_MAX_FAWC_P1_S6
`endif 

`ifdef i_axi_AXI_MAX_FARC_S6
  `define AXI_MAX_FARC_S6 `i_axi_AXI_MAX_FARC_S6
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FARC_P1_S6
  `define AXI_LOG2_MAX_FARC_P1_S6 `i_axi_AXI_LOG2_MAX_FARC_P1_S6
`endif 

`ifdef i_axi_AXI_WID_S7
  `define AXI_WID_S7 `i_axi_AXI_WID_S7
`endif 

`ifdef i_axi_AXI_LOG2_WID_S7
  `define AXI_LOG2_WID_S7 `i_axi_AXI_LOG2_WID_S7
`endif 

`ifdef i_axi_AXI_LOG2_WID_P1_S7
  `define AXI_LOG2_WID_P1_S7 `i_axi_AXI_LOG2_WID_P1_S7
`endif 

`ifdef i_axi_AXI_MAX_FAWC_S7
  `define AXI_MAX_FAWC_S7 `i_axi_AXI_MAX_FAWC_S7
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_S7
  `define AXI_LOG2_MAX_FAWC_S7 `i_axi_AXI_LOG2_MAX_FAWC_S7
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_P1_S7
  `define AXI_LOG2_MAX_FAWC_P1_S7 `i_axi_AXI_LOG2_MAX_FAWC_P1_S7
`endif 

`ifdef i_axi_AXI_MAX_FARC_S7
  `define AXI_MAX_FARC_S7 `i_axi_AXI_MAX_FARC_S7
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FARC_P1_S7
  `define AXI_LOG2_MAX_FARC_P1_S7 `i_axi_AXI_LOG2_MAX_FARC_P1_S7
`endif 

`ifdef i_axi_AXI_WID_S8
  `define AXI_WID_S8 `i_axi_AXI_WID_S8
`endif 

`ifdef i_axi_AXI_LOG2_WID_S8
  `define AXI_LOG2_WID_S8 `i_axi_AXI_LOG2_WID_S8
`endif 

`ifdef i_axi_AXI_LOG2_WID_P1_S8
  `define AXI_LOG2_WID_P1_S8 `i_axi_AXI_LOG2_WID_P1_S8
`endif 

`ifdef i_axi_AXI_MAX_FAWC_S8
  `define AXI_MAX_FAWC_S8 `i_axi_AXI_MAX_FAWC_S8
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_S8
  `define AXI_LOG2_MAX_FAWC_S8 `i_axi_AXI_LOG2_MAX_FAWC_S8
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_P1_S8
  `define AXI_LOG2_MAX_FAWC_P1_S8 `i_axi_AXI_LOG2_MAX_FAWC_P1_S8
`endif 

`ifdef i_axi_AXI_MAX_FARC_S8
  `define AXI_MAX_FARC_S8 `i_axi_AXI_MAX_FARC_S8
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FARC_P1_S8
  `define AXI_LOG2_MAX_FARC_P1_S8 `i_axi_AXI_LOG2_MAX_FARC_P1_S8
`endif 

`ifdef i_axi_AXI_WID_S9
  `define AXI_WID_S9 `i_axi_AXI_WID_S9
`endif 

`ifdef i_axi_AXI_LOG2_WID_S9
  `define AXI_LOG2_WID_S9 `i_axi_AXI_LOG2_WID_S9
`endif 

`ifdef i_axi_AXI_LOG2_WID_P1_S9
  `define AXI_LOG2_WID_P1_S9 `i_axi_AXI_LOG2_WID_P1_S9
`endif 

`ifdef i_axi_AXI_MAX_FAWC_S9
  `define AXI_MAX_FAWC_S9 `i_axi_AXI_MAX_FAWC_S9
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_S9
  `define AXI_LOG2_MAX_FAWC_S9 `i_axi_AXI_LOG2_MAX_FAWC_S9
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_P1_S9
  `define AXI_LOG2_MAX_FAWC_P1_S9 `i_axi_AXI_LOG2_MAX_FAWC_P1_S9
`endif 

`ifdef i_axi_AXI_MAX_FARC_S9
  `define AXI_MAX_FARC_S9 `i_axi_AXI_MAX_FARC_S9
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FARC_P1_S9
  `define AXI_LOG2_MAX_FARC_P1_S9 `i_axi_AXI_LOG2_MAX_FARC_P1_S9
`endif 

`ifdef i_axi_AXI_WID_S10
  `define AXI_WID_S10 `i_axi_AXI_WID_S10
`endif 

`ifdef i_axi_AXI_LOG2_WID_S10
  `define AXI_LOG2_WID_S10 `i_axi_AXI_LOG2_WID_S10
`endif 

`ifdef i_axi_AXI_LOG2_WID_P1_S10
  `define AXI_LOG2_WID_P1_S10 `i_axi_AXI_LOG2_WID_P1_S10
`endif 

`ifdef i_axi_AXI_MAX_FAWC_S10
  `define AXI_MAX_FAWC_S10 `i_axi_AXI_MAX_FAWC_S10
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_S10
  `define AXI_LOG2_MAX_FAWC_S10 `i_axi_AXI_LOG2_MAX_FAWC_S10
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_P1_S10
  `define AXI_LOG2_MAX_FAWC_P1_S10 `i_axi_AXI_LOG2_MAX_FAWC_P1_S10
`endif 

`ifdef i_axi_AXI_MAX_FARC_S10
  `define AXI_MAX_FARC_S10 `i_axi_AXI_MAX_FARC_S10
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FARC_P1_S10
  `define AXI_LOG2_MAX_FARC_P1_S10 `i_axi_AXI_LOG2_MAX_FARC_P1_S10
`endif 

`ifdef i_axi_AXI_WID_S11
  `define AXI_WID_S11 `i_axi_AXI_WID_S11
`endif 

`ifdef i_axi_AXI_LOG2_WID_S11
  `define AXI_LOG2_WID_S11 `i_axi_AXI_LOG2_WID_S11
`endif 

`ifdef i_axi_AXI_LOG2_WID_P1_S11
  `define AXI_LOG2_WID_P1_S11 `i_axi_AXI_LOG2_WID_P1_S11
`endif 

`ifdef i_axi_AXI_MAX_FAWC_S11
  `define AXI_MAX_FAWC_S11 `i_axi_AXI_MAX_FAWC_S11
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_S11
  `define AXI_LOG2_MAX_FAWC_S11 `i_axi_AXI_LOG2_MAX_FAWC_S11
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_P1_S11
  `define AXI_LOG2_MAX_FAWC_P1_S11 `i_axi_AXI_LOG2_MAX_FAWC_P1_S11
`endif 

`ifdef i_axi_AXI_MAX_FARC_S11
  `define AXI_MAX_FARC_S11 `i_axi_AXI_MAX_FARC_S11
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FARC_P1_S11
  `define AXI_LOG2_MAX_FARC_P1_S11 `i_axi_AXI_LOG2_MAX_FARC_P1_S11
`endif 

`ifdef i_axi_AXI_WID_S12
  `define AXI_WID_S12 `i_axi_AXI_WID_S12
`endif 

`ifdef i_axi_AXI_LOG2_WID_S12
  `define AXI_LOG2_WID_S12 `i_axi_AXI_LOG2_WID_S12
`endif 

`ifdef i_axi_AXI_LOG2_WID_P1_S12
  `define AXI_LOG2_WID_P1_S12 `i_axi_AXI_LOG2_WID_P1_S12
`endif 

`ifdef i_axi_AXI_MAX_FAWC_S12
  `define AXI_MAX_FAWC_S12 `i_axi_AXI_MAX_FAWC_S12
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_S12
  `define AXI_LOG2_MAX_FAWC_S12 `i_axi_AXI_LOG2_MAX_FAWC_S12
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_P1_S12
  `define AXI_LOG2_MAX_FAWC_P1_S12 `i_axi_AXI_LOG2_MAX_FAWC_P1_S12
`endif 

`ifdef i_axi_AXI_MAX_FARC_S12
  `define AXI_MAX_FARC_S12 `i_axi_AXI_MAX_FARC_S12
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FARC_P1_S12
  `define AXI_LOG2_MAX_FARC_P1_S12 `i_axi_AXI_LOG2_MAX_FARC_P1_S12
`endif 

`ifdef i_axi_AXI_WID_S13
  `define AXI_WID_S13 `i_axi_AXI_WID_S13
`endif 

`ifdef i_axi_AXI_LOG2_WID_S13
  `define AXI_LOG2_WID_S13 `i_axi_AXI_LOG2_WID_S13
`endif 

`ifdef i_axi_AXI_LOG2_WID_P1_S13
  `define AXI_LOG2_WID_P1_S13 `i_axi_AXI_LOG2_WID_P1_S13
`endif 

`ifdef i_axi_AXI_MAX_FAWC_S13
  `define AXI_MAX_FAWC_S13 `i_axi_AXI_MAX_FAWC_S13
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_S13
  `define AXI_LOG2_MAX_FAWC_S13 `i_axi_AXI_LOG2_MAX_FAWC_S13
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_P1_S13
  `define AXI_LOG2_MAX_FAWC_P1_S13 `i_axi_AXI_LOG2_MAX_FAWC_P1_S13
`endif 

`ifdef i_axi_AXI_MAX_FARC_S13
  `define AXI_MAX_FARC_S13 `i_axi_AXI_MAX_FARC_S13
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FARC_P1_S13
  `define AXI_LOG2_MAX_FARC_P1_S13 `i_axi_AXI_LOG2_MAX_FARC_P1_S13
`endif 

`ifdef i_axi_AXI_WID_S14
  `define AXI_WID_S14 `i_axi_AXI_WID_S14
`endif 

`ifdef i_axi_AXI_LOG2_WID_S14
  `define AXI_LOG2_WID_S14 `i_axi_AXI_LOG2_WID_S14
`endif 

`ifdef i_axi_AXI_LOG2_WID_P1_S14
  `define AXI_LOG2_WID_P1_S14 `i_axi_AXI_LOG2_WID_P1_S14
`endif 

`ifdef i_axi_AXI_MAX_FAWC_S14
  `define AXI_MAX_FAWC_S14 `i_axi_AXI_MAX_FAWC_S14
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_S14
  `define AXI_LOG2_MAX_FAWC_S14 `i_axi_AXI_LOG2_MAX_FAWC_S14
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_P1_S14
  `define AXI_LOG2_MAX_FAWC_P1_S14 `i_axi_AXI_LOG2_MAX_FAWC_P1_S14
`endif 

`ifdef i_axi_AXI_MAX_FARC_S14
  `define AXI_MAX_FARC_S14 `i_axi_AXI_MAX_FARC_S14
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FARC_P1_S14
  `define AXI_LOG2_MAX_FARC_P1_S14 `i_axi_AXI_LOG2_MAX_FARC_P1_S14
`endif 

`ifdef i_axi_AXI_WID_S15
  `define AXI_WID_S15 `i_axi_AXI_WID_S15
`endif 

`ifdef i_axi_AXI_LOG2_WID_S15
  `define AXI_LOG2_WID_S15 `i_axi_AXI_LOG2_WID_S15
`endif 

`ifdef i_axi_AXI_LOG2_WID_P1_S15
  `define AXI_LOG2_WID_P1_S15 `i_axi_AXI_LOG2_WID_P1_S15
`endif 

`ifdef i_axi_AXI_MAX_FAWC_S15
  `define AXI_MAX_FAWC_S15 `i_axi_AXI_MAX_FAWC_S15
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_S15
  `define AXI_LOG2_MAX_FAWC_S15 `i_axi_AXI_LOG2_MAX_FAWC_S15
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_P1_S15
  `define AXI_LOG2_MAX_FAWC_P1_S15 `i_axi_AXI_LOG2_MAX_FAWC_P1_S15
`endif 

`ifdef i_axi_AXI_MAX_FARC_S15
  `define AXI_MAX_FARC_S15 `i_axi_AXI_MAX_FARC_S15
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FARC_P1_S15
  `define AXI_LOG2_MAX_FARC_P1_S15 `i_axi_AXI_LOG2_MAX_FARC_P1_S15
`endif 

`ifdef i_axi_AXI_WID_S16
  `define AXI_WID_S16 `i_axi_AXI_WID_S16
`endif 

`ifdef i_axi_AXI_LOG2_WID_S16
  `define AXI_LOG2_WID_S16 `i_axi_AXI_LOG2_WID_S16
`endif 

`ifdef i_axi_AXI_LOG2_WID_P1_S16
  `define AXI_LOG2_WID_P1_S16 `i_axi_AXI_LOG2_WID_P1_S16
`endif 

`ifdef i_axi_AXI_MAX_FAWC_S16
  `define AXI_MAX_FAWC_S16 `i_axi_AXI_MAX_FAWC_S16
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_S16
  `define AXI_LOG2_MAX_FAWC_S16 `i_axi_AXI_LOG2_MAX_FAWC_S16
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FAWC_P1_S16
  `define AXI_LOG2_MAX_FAWC_P1_S16 `i_axi_AXI_LOG2_MAX_FAWC_P1_S16
`endif 

`ifdef i_axi_AXI_MAX_FARC_S16
  `define AXI_MAX_FARC_S16 `i_axi_AXI_MAX_FARC_S16
`endif 

`ifdef i_axi_AXI_LOG2_MAX_FARC_P1_S16
  `define AXI_LOG2_MAX_FARC_P1_S16 `i_axi_AXI_LOG2_MAX_FARC_P1_S16
`endif 

`ifdef i_axi_AXI_S0_SHARED_FARC
  `define AXI_S0_SHARED_FARC `i_axi_AXI_S0_SHARED_FARC
`endif 

`ifdef i_axi_AXI_LOG2_S0_SHARED_FARC_P1
  `define AXI_LOG2_S0_SHARED_FARC_P1 `i_axi_AXI_LOG2_S0_SHARED_FARC_P1
`endif 

`ifdef i_axi_AXI_S0_SHARED_AR_HAS_DDCTD
  `define AXI_S0_SHARED_AR_HAS_DDCTD `i_axi_AXI_S0_SHARED_AR_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S0_SHARED_FAWC
  `define AXI_S0_SHARED_FAWC `i_axi_AXI_S0_SHARED_FAWC
`endif 

`ifdef i_axi_AXI_LOG2_S0_SHARED_FAWC_P1
  `define AXI_LOG2_S0_SHARED_FAWC_P1 `i_axi_AXI_LOG2_S0_SHARED_FAWC_P1
`endif 

`ifdef i_axi_AXI_S0_SHARED_AW_HAS_DDCTD
  `define AXI_S0_SHARED_AW_HAS_DDCTD `i_axi_AXI_S0_SHARED_AW_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S0_SHARED_W_HAS_DDCTD
  `define AXI_S0_SHARED_W_HAS_DDCTD `i_axi_AXI_S0_SHARED_W_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S1_SHARED_FARC
  `define AXI_S1_SHARED_FARC `i_axi_AXI_S1_SHARED_FARC
`endif 

`ifdef i_axi_AXI_LOG2_S1_SHARED_FARC_P1
  `define AXI_LOG2_S1_SHARED_FARC_P1 `i_axi_AXI_LOG2_S1_SHARED_FARC_P1
`endif 

`ifdef i_axi_AXI_S1_SHARED_AR_HAS_DDCTD
  `define AXI_S1_SHARED_AR_HAS_DDCTD `i_axi_AXI_S1_SHARED_AR_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S1_SHARED_FAWC
  `define AXI_S1_SHARED_FAWC `i_axi_AXI_S1_SHARED_FAWC
`endif 

`ifdef i_axi_AXI_LOG2_S1_SHARED_FAWC_P1
  `define AXI_LOG2_S1_SHARED_FAWC_P1 `i_axi_AXI_LOG2_S1_SHARED_FAWC_P1
`endif 

`ifdef i_axi_AXI_S1_SHARED_AW_HAS_DDCTD
  `define AXI_S1_SHARED_AW_HAS_DDCTD `i_axi_AXI_S1_SHARED_AW_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S1_SHARED_W_HAS_DDCTD
  `define AXI_S1_SHARED_W_HAS_DDCTD `i_axi_AXI_S1_SHARED_W_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S2_SHARED_FARC
  `define AXI_S2_SHARED_FARC `i_axi_AXI_S2_SHARED_FARC
`endif 

`ifdef i_axi_AXI_LOG2_S2_SHARED_FARC_P1
  `define AXI_LOG2_S2_SHARED_FARC_P1 `i_axi_AXI_LOG2_S2_SHARED_FARC_P1
`endif 

`ifdef i_axi_AXI_S2_SHARED_AR_HAS_DDCTD
  `define AXI_S2_SHARED_AR_HAS_DDCTD `i_axi_AXI_S2_SHARED_AR_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S2_SHARED_FAWC
  `define AXI_S2_SHARED_FAWC `i_axi_AXI_S2_SHARED_FAWC
`endif 

`ifdef i_axi_AXI_LOG2_S2_SHARED_FAWC_P1
  `define AXI_LOG2_S2_SHARED_FAWC_P1 `i_axi_AXI_LOG2_S2_SHARED_FAWC_P1
`endif 

`ifdef i_axi_AXI_S2_SHARED_AW_HAS_DDCTD
  `define AXI_S2_SHARED_AW_HAS_DDCTD `i_axi_AXI_S2_SHARED_AW_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S2_SHARED_W_HAS_DDCTD
  `define AXI_S2_SHARED_W_HAS_DDCTD `i_axi_AXI_S2_SHARED_W_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S3_SHARED_FARC
  `define AXI_S3_SHARED_FARC `i_axi_AXI_S3_SHARED_FARC
`endif 

`ifdef i_axi_AXI_LOG2_S3_SHARED_FARC_P1
  `define AXI_LOG2_S3_SHARED_FARC_P1 `i_axi_AXI_LOG2_S3_SHARED_FARC_P1
`endif 

`ifdef i_axi_AXI_S3_SHARED_AR_HAS_DDCTD
  `define AXI_S3_SHARED_AR_HAS_DDCTD `i_axi_AXI_S3_SHARED_AR_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S3_SHARED_FAWC
  `define AXI_S3_SHARED_FAWC `i_axi_AXI_S3_SHARED_FAWC
`endif 

`ifdef i_axi_AXI_LOG2_S3_SHARED_FAWC_P1
  `define AXI_LOG2_S3_SHARED_FAWC_P1 `i_axi_AXI_LOG2_S3_SHARED_FAWC_P1
`endif 

`ifdef i_axi_AXI_S3_SHARED_AW_HAS_DDCTD
  `define AXI_S3_SHARED_AW_HAS_DDCTD `i_axi_AXI_S3_SHARED_AW_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S3_SHARED_W_HAS_DDCTD
  `define AXI_S3_SHARED_W_HAS_DDCTD `i_axi_AXI_S3_SHARED_W_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S4_SHARED_FARC
  `define AXI_S4_SHARED_FARC `i_axi_AXI_S4_SHARED_FARC
`endif 

`ifdef i_axi_AXI_LOG2_S4_SHARED_FARC_P1
  `define AXI_LOG2_S4_SHARED_FARC_P1 `i_axi_AXI_LOG2_S4_SHARED_FARC_P1
`endif 

`ifdef i_axi_AXI_S4_SHARED_AR_HAS_DDCTD
  `define AXI_S4_SHARED_AR_HAS_DDCTD `i_axi_AXI_S4_SHARED_AR_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S4_SHARED_FAWC
  `define AXI_S4_SHARED_FAWC `i_axi_AXI_S4_SHARED_FAWC
`endif 

`ifdef i_axi_AXI_LOG2_S4_SHARED_FAWC_P1
  `define AXI_LOG2_S4_SHARED_FAWC_P1 `i_axi_AXI_LOG2_S4_SHARED_FAWC_P1
`endif 

`ifdef i_axi_AXI_S4_SHARED_AW_HAS_DDCTD
  `define AXI_S4_SHARED_AW_HAS_DDCTD `i_axi_AXI_S4_SHARED_AW_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S4_SHARED_W_HAS_DDCTD
  `define AXI_S4_SHARED_W_HAS_DDCTD `i_axi_AXI_S4_SHARED_W_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S5_SHARED_FARC
  `define AXI_S5_SHARED_FARC `i_axi_AXI_S5_SHARED_FARC
`endif 

`ifdef i_axi_AXI_LOG2_S5_SHARED_FARC_P1
  `define AXI_LOG2_S5_SHARED_FARC_P1 `i_axi_AXI_LOG2_S5_SHARED_FARC_P1
`endif 

`ifdef i_axi_AXI_S5_SHARED_AR_HAS_DDCTD
  `define AXI_S5_SHARED_AR_HAS_DDCTD `i_axi_AXI_S5_SHARED_AR_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S5_SHARED_FAWC
  `define AXI_S5_SHARED_FAWC `i_axi_AXI_S5_SHARED_FAWC
`endif 

`ifdef i_axi_AXI_LOG2_S5_SHARED_FAWC_P1
  `define AXI_LOG2_S5_SHARED_FAWC_P1 `i_axi_AXI_LOG2_S5_SHARED_FAWC_P1
`endif 

`ifdef i_axi_AXI_S5_SHARED_AW_HAS_DDCTD
  `define AXI_S5_SHARED_AW_HAS_DDCTD `i_axi_AXI_S5_SHARED_AW_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S5_SHARED_W_HAS_DDCTD
  `define AXI_S5_SHARED_W_HAS_DDCTD `i_axi_AXI_S5_SHARED_W_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S6_SHARED_FARC
  `define AXI_S6_SHARED_FARC `i_axi_AXI_S6_SHARED_FARC
`endif 

`ifdef i_axi_AXI_LOG2_S6_SHARED_FARC_P1
  `define AXI_LOG2_S6_SHARED_FARC_P1 `i_axi_AXI_LOG2_S6_SHARED_FARC_P1
`endif 

`ifdef i_axi_AXI_S6_SHARED_AR_HAS_DDCTD
  `define AXI_S6_SHARED_AR_HAS_DDCTD `i_axi_AXI_S6_SHARED_AR_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S6_SHARED_FAWC
  `define AXI_S6_SHARED_FAWC `i_axi_AXI_S6_SHARED_FAWC
`endif 

`ifdef i_axi_AXI_LOG2_S6_SHARED_FAWC_P1
  `define AXI_LOG2_S6_SHARED_FAWC_P1 `i_axi_AXI_LOG2_S6_SHARED_FAWC_P1
`endif 

`ifdef i_axi_AXI_S6_SHARED_AW_HAS_DDCTD
  `define AXI_S6_SHARED_AW_HAS_DDCTD `i_axi_AXI_S6_SHARED_AW_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S6_SHARED_W_HAS_DDCTD
  `define AXI_S6_SHARED_W_HAS_DDCTD `i_axi_AXI_S6_SHARED_W_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S7_SHARED_FARC
  `define AXI_S7_SHARED_FARC `i_axi_AXI_S7_SHARED_FARC
`endif 

`ifdef i_axi_AXI_LOG2_S7_SHARED_FARC_P1
  `define AXI_LOG2_S7_SHARED_FARC_P1 `i_axi_AXI_LOG2_S7_SHARED_FARC_P1
`endif 

`ifdef i_axi_AXI_S7_SHARED_AR_HAS_DDCTD
  `define AXI_S7_SHARED_AR_HAS_DDCTD `i_axi_AXI_S7_SHARED_AR_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S7_SHARED_FAWC
  `define AXI_S7_SHARED_FAWC `i_axi_AXI_S7_SHARED_FAWC
`endif 

`ifdef i_axi_AXI_LOG2_S7_SHARED_FAWC_P1
  `define AXI_LOG2_S7_SHARED_FAWC_P1 `i_axi_AXI_LOG2_S7_SHARED_FAWC_P1
`endif 

`ifdef i_axi_AXI_S7_SHARED_AW_HAS_DDCTD
  `define AXI_S7_SHARED_AW_HAS_DDCTD `i_axi_AXI_S7_SHARED_AW_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S7_SHARED_W_HAS_DDCTD
  `define AXI_S7_SHARED_W_HAS_DDCTD `i_axi_AXI_S7_SHARED_W_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S8_SHARED_FARC
  `define AXI_S8_SHARED_FARC `i_axi_AXI_S8_SHARED_FARC
`endif 

`ifdef i_axi_AXI_LOG2_S8_SHARED_FARC_P1
  `define AXI_LOG2_S8_SHARED_FARC_P1 `i_axi_AXI_LOG2_S8_SHARED_FARC_P1
`endif 

`ifdef i_axi_AXI_S8_SHARED_AR_HAS_DDCTD
  `define AXI_S8_SHARED_AR_HAS_DDCTD `i_axi_AXI_S8_SHARED_AR_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S8_SHARED_FAWC
  `define AXI_S8_SHARED_FAWC `i_axi_AXI_S8_SHARED_FAWC
`endif 

`ifdef i_axi_AXI_LOG2_S8_SHARED_FAWC_P1
  `define AXI_LOG2_S8_SHARED_FAWC_P1 `i_axi_AXI_LOG2_S8_SHARED_FAWC_P1
`endif 

`ifdef i_axi_AXI_S8_SHARED_AW_HAS_DDCTD
  `define AXI_S8_SHARED_AW_HAS_DDCTD `i_axi_AXI_S8_SHARED_AW_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S8_SHARED_W_HAS_DDCTD
  `define AXI_S8_SHARED_W_HAS_DDCTD `i_axi_AXI_S8_SHARED_W_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S9_SHARED_FARC
  `define AXI_S9_SHARED_FARC `i_axi_AXI_S9_SHARED_FARC
`endif 

`ifdef i_axi_AXI_LOG2_S9_SHARED_FARC_P1
  `define AXI_LOG2_S9_SHARED_FARC_P1 `i_axi_AXI_LOG2_S9_SHARED_FARC_P1
`endif 

`ifdef i_axi_AXI_S9_SHARED_AR_HAS_DDCTD
  `define AXI_S9_SHARED_AR_HAS_DDCTD `i_axi_AXI_S9_SHARED_AR_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S9_SHARED_FAWC
  `define AXI_S9_SHARED_FAWC `i_axi_AXI_S9_SHARED_FAWC
`endif 

`ifdef i_axi_AXI_LOG2_S9_SHARED_FAWC_P1
  `define AXI_LOG2_S9_SHARED_FAWC_P1 `i_axi_AXI_LOG2_S9_SHARED_FAWC_P1
`endif 

`ifdef i_axi_AXI_S9_SHARED_AW_HAS_DDCTD
  `define AXI_S9_SHARED_AW_HAS_DDCTD `i_axi_AXI_S9_SHARED_AW_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S9_SHARED_W_HAS_DDCTD
  `define AXI_S9_SHARED_W_HAS_DDCTD `i_axi_AXI_S9_SHARED_W_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S10_SHARED_FARC
  `define AXI_S10_SHARED_FARC `i_axi_AXI_S10_SHARED_FARC
`endif 

`ifdef i_axi_AXI_LOG2_S10_SHARED_FARC_P1
  `define AXI_LOG2_S10_SHARED_FARC_P1 `i_axi_AXI_LOG2_S10_SHARED_FARC_P1
`endif 

`ifdef i_axi_AXI_S10_SHARED_AR_HAS_DDCTD
  `define AXI_S10_SHARED_AR_HAS_DDCTD `i_axi_AXI_S10_SHARED_AR_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S10_SHARED_FAWC
  `define AXI_S10_SHARED_FAWC `i_axi_AXI_S10_SHARED_FAWC
`endif 

`ifdef i_axi_AXI_LOG2_S10_SHARED_FAWC_P1
  `define AXI_LOG2_S10_SHARED_FAWC_P1 `i_axi_AXI_LOG2_S10_SHARED_FAWC_P1
`endif 

`ifdef i_axi_AXI_S10_SHARED_AW_HAS_DDCTD
  `define AXI_S10_SHARED_AW_HAS_DDCTD `i_axi_AXI_S10_SHARED_AW_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S10_SHARED_W_HAS_DDCTD
  `define AXI_S10_SHARED_W_HAS_DDCTD `i_axi_AXI_S10_SHARED_W_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S11_SHARED_FARC
  `define AXI_S11_SHARED_FARC `i_axi_AXI_S11_SHARED_FARC
`endif 

`ifdef i_axi_AXI_LOG2_S11_SHARED_FARC_P1
  `define AXI_LOG2_S11_SHARED_FARC_P1 `i_axi_AXI_LOG2_S11_SHARED_FARC_P1
`endif 

`ifdef i_axi_AXI_S11_SHARED_AR_HAS_DDCTD
  `define AXI_S11_SHARED_AR_HAS_DDCTD `i_axi_AXI_S11_SHARED_AR_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S11_SHARED_FAWC
  `define AXI_S11_SHARED_FAWC `i_axi_AXI_S11_SHARED_FAWC
`endif 

`ifdef i_axi_AXI_LOG2_S11_SHARED_FAWC_P1
  `define AXI_LOG2_S11_SHARED_FAWC_P1 `i_axi_AXI_LOG2_S11_SHARED_FAWC_P1
`endif 

`ifdef i_axi_AXI_S11_SHARED_AW_HAS_DDCTD
  `define AXI_S11_SHARED_AW_HAS_DDCTD `i_axi_AXI_S11_SHARED_AW_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S11_SHARED_W_HAS_DDCTD
  `define AXI_S11_SHARED_W_HAS_DDCTD `i_axi_AXI_S11_SHARED_W_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S12_SHARED_FARC
  `define AXI_S12_SHARED_FARC `i_axi_AXI_S12_SHARED_FARC
`endif 

`ifdef i_axi_AXI_LOG2_S12_SHARED_FARC_P1
  `define AXI_LOG2_S12_SHARED_FARC_P1 `i_axi_AXI_LOG2_S12_SHARED_FARC_P1
`endif 

`ifdef i_axi_AXI_S12_SHARED_AR_HAS_DDCTD
  `define AXI_S12_SHARED_AR_HAS_DDCTD `i_axi_AXI_S12_SHARED_AR_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S12_SHARED_FAWC
  `define AXI_S12_SHARED_FAWC `i_axi_AXI_S12_SHARED_FAWC
`endif 

`ifdef i_axi_AXI_LOG2_S12_SHARED_FAWC_P1
  `define AXI_LOG2_S12_SHARED_FAWC_P1 `i_axi_AXI_LOG2_S12_SHARED_FAWC_P1
`endif 

`ifdef i_axi_AXI_S12_SHARED_AW_HAS_DDCTD
  `define AXI_S12_SHARED_AW_HAS_DDCTD `i_axi_AXI_S12_SHARED_AW_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S12_SHARED_W_HAS_DDCTD
  `define AXI_S12_SHARED_W_HAS_DDCTD `i_axi_AXI_S12_SHARED_W_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S13_SHARED_FARC
  `define AXI_S13_SHARED_FARC `i_axi_AXI_S13_SHARED_FARC
`endif 

`ifdef i_axi_AXI_LOG2_S13_SHARED_FARC_P1
  `define AXI_LOG2_S13_SHARED_FARC_P1 `i_axi_AXI_LOG2_S13_SHARED_FARC_P1
`endif 

`ifdef i_axi_AXI_S13_SHARED_AR_HAS_DDCTD
  `define AXI_S13_SHARED_AR_HAS_DDCTD `i_axi_AXI_S13_SHARED_AR_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S13_SHARED_FAWC
  `define AXI_S13_SHARED_FAWC `i_axi_AXI_S13_SHARED_FAWC
`endif 

`ifdef i_axi_AXI_LOG2_S13_SHARED_FAWC_P1
  `define AXI_LOG2_S13_SHARED_FAWC_P1 `i_axi_AXI_LOG2_S13_SHARED_FAWC_P1
`endif 

`ifdef i_axi_AXI_S13_SHARED_AW_HAS_DDCTD
  `define AXI_S13_SHARED_AW_HAS_DDCTD `i_axi_AXI_S13_SHARED_AW_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S13_SHARED_W_HAS_DDCTD
  `define AXI_S13_SHARED_W_HAS_DDCTD `i_axi_AXI_S13_SHARED_W_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S14_SHARED_FARC
  `define AXI_S14_SHARED_FARC `i_axi_AXI_S14_SHARED_FARC
`endif 

`ifdef i_axi_AXI_LOG2_S14_SHARED_FARC_P1
  `define AXI_LOG2_S14_SHARED_FARC_P1 `i_axi_AXI_LOG2_S14_SHARED_FARC_P1
`endif 

`ifdef i_axi_AXI_S14_SHARED_AR_HAS_DDCTD
  `define AXI_S14_SHARED_AR_HAS_DDCTD `i_axi_AXI_S14_SHARED_AR_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S14_SHARED_FAWC
  `define AXI_S14_SHARED_FAWC `i_axi_AXI_S14_SHARED_FAWC
`endif 

`ifdef i_axi_AXI_LOG2_S14_SHARED_FAWC_P1
  `define AXI_LOG2_S14_SHARED_FAWC_P1 `i_axi_AXI_LOG2_S14_SHARED_FAWC_P1
`endif 

`ifdef i_axi_AXI_S14_SHARED_AW_HAS_DDCTD
  `define AXI_S14_SHARED_AW_HAS_DDCTD `i_axi_AXI_S14_SHARED_AW_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S14_SHARED_W_HAS_DDCTD
  `define AXI_S14_SHARED_W_HAS_DDCTD `i_axi_AXI_S14_SHARED_W_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S15_SHARED_FARC
  `define AXI_S15_SHARED_FARC `i_axi_AXI_S15_SHARED_FARC
`endif 

`ifdef i_axi_AXI_LOG2_S15_SHARED_FARC_P1
  `define AXI_LOG2_S15_SHARED_FARC_P1 `i_axi_AXI_LOG2_S15_SHARED_FARC_P1
`endif 

`ifdef i_axi_AXI_S15_SHARED_AR_HAS_DDCTD
  `define AXI_S15_SHARED_AR_HAS_DDCTD `i_axi_AXI_S15_SHARED_AR_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S15_SHARED_FAWC
  `define AXI_S15_SHARED_FAWC `i_axi_AXI_S15_SHARED_FAWC
`endif 

`ifdef i_axi_AXI_LOG2_S15_SHARED_FAWC_P1
  `define AXI_LOG2_S15_SHARED_FAWC_P1 `i_axi_AXI_LOG2_S15_SHARED_FAWC_P1
`endif 

`ifdef i_axi_AXI_S15_SHARED_AW_HAS_DDCTD
  `define AXI_S15_SHARED_AW_HAS_DDCTD `i_axi_AXI_S15_SHARED_AW_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S15_SHARED_W_HAS_DDCTD
  `define AXI_S15_SHARED_W_HAS_DDCTD `i_axi_AXI_S15_SHARED_W_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S16_SHARED_FARC
  `define AXI_S16_SHARED_FARC `i_axi_AXI_S16_SHARED_FARC
`endif 

`ifdef i_axi_AXI_LOG2_S16_SHARED_FARC_P1
  `define AXI_LOG2_S16_SHARED_FARC_P1 `i_axi_AXI_LOG2_S16_SHARED_FARC_P1
`endif 

`ifdef i_axi_AXI_S16_SHARED_AR_HAS_DDCTD
  `define AXI_S16_SHARED_AR_HAS_DDCTD `i_axi_AXI_S16_SHARED_AR_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S16_SHARED_FAWC
  `define AXI_S16_SHARED_FAWC `i_axi_AXI_S16_SHARED_FAWC
`endif 

`ifdef i_axi_AXI_LOG2_S16_SHARED_FAWC_P1
  `define AXI_LOG2_S16_SHARED_FAWC_P1 `i_axi_AXI_LOG2_S16_SHARED_FAWC_P1
`endif 

`ifdef i_axi_AXI_S16_SHARED_AW_HAS_DDCTD
  `define AXI_S16_SHARED_AW_HAS_DDCTD `i_axi_AXI_S16_SHARED_AW_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_S16_SHARED_W_HAS_DDCTD
  `define AXI_S16_SHARED_W_HAS_DDCTD `i_axi_AXI_S16_SHARED_W_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M0_SHARED_R_HAS_DDCTD
  `define AXI_M0_SHARED_R_HAS_DDCTD `i_axi_AXI_M0_SHARED_R_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M0_SHARED_B_HAS_DDCTD
  `define AXI_M0_SHARED_B_HAS_DDCTD `i_axi_AXI_M0_SHARED_B_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M1_SHARED_R_HAS_DDCTD
  `define AXI_M1_SHARED_R_HAS_DDCTD `i_axi_AXI_M1_SHARED_R_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M1_SHARED_B_HAS_DDCTD
  `define AXI_M1_SHARED_B_HAS_DDCTD `i_axi_AXI_M1_SHARED_B_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M2_SHARED_R_HAS_DDCTD
  `define AXI_M2_SHARED_R_HAS_DDCTD `i_axi_AXI_M2_SHARED_R_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M2_SHARED_B_HAS_DDCTD
  `define AXI_M2_SHARED_B_HAS_DDCTD `i_axi_AXI_M2_SHARED_B_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M3_SHARED_R_HAS_DDCTD
  `define AXI_M3_SHARED_R_HAS_DDCTD `i_axi_AXI_M3_SHARED_R_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M3_SHARED_B_HAS_DDCTD
  `define AXI_M3_SHARED_B_HAS_DDCTD `i_axi_AXI_M3_SHARED_B_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M4_SHARED_R_HAS_DDCTD
  `define AXI_M4_SHARED_R_HAS_DDCTD `i_axi_AXI_M4_SHARED_R_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M4_SHARED_B_HAS_DDCTD
  `define AXI_M4_SHARED_B_HAS_DDCTD `i_axi_AXI_M4_SHARED_B_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M5_SHARED_R_HAS_DDCTD
  `define AXI_M5_SHARED_R_HAS_DDCTD `i_axi_AXI_M5_SHARED_R_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M5_SHARED_B_HAS_DDCTD
  `define AXI_M5_SHARED_B_HAS_DDCTD `i_axi_AXI_M5_SHARED_B_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M6_SHARED_R_HAS_DDCTD
  `define AXI_M6_SHARED_R_HAS_DDCTD `i_axi_AXI_M6_SHARED_R_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M6_SHARED_B_HAS_DDCTD
  `define AXI_M6_SHARED_B_HAS_DDCTD `i_axi_AXI_M6_SHARED_B_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M7_SHARED_R_HAS_DDCTD
  `define AXI_M7_SHARED_R_HAS_DDCTD `i_axi_AXI_M7_SHARED_R_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M7_SHARED_B_HAS_DDCTD
  `define AXI_M7_SHARED_B_HAS_DDCTD `i_axi_AXI_M7_SHARED_B_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M8_SHARED_R_HAS_DDCTD
  `define AXI_M8_SHARED_R_HAS_DDCTD `i_axi_AXI_M8_SHARED_R_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M8_SHARED_B_HAS_DDCTD
  `define AXI_M8_SHARED_B_HAS_DDCTD `i_axi_AXI_M8_SHARED_B_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M9_SHARED_R_HAS_DDCTD
  `define AXI_M9_SHARED_R_HAS_DDCTD `i_axi_AXI_M9_SHARED_R_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M9_SHARED_B_HAS_DDCTD
  `define AXI_M9_SHARED_B_HAS_DDCTD `i_axi_AXI_M9_SHARED_B_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M10_SHARED_R_HAS_DDCTD
  `define AXI_M10_SHARED_R_HAS_DDCTD `i_axi_AXI_M10_SHARED_R_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M10_SHARED_B_HAS_DDCTD
  `define AXI_M10_SHARED_B_HAS_DDCTD `i_axi_AXI_M10_SHARED_B_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M11_SHARED_R_HAS_DDCTD
  `define AXI_M11_SHARED_R_HAS_DDCTD `i_axi_AXI_M11_SHARED_R_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M11_SHARED_B_HAS_DDCTD
  `define AXI_M11_SHARED_B_HAS_DDCTD `i_axi_AXI_M11_SHARED_B_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M12_SHARED_R_HAS_DDCTD
  `define AXI_M12_SHARED_R_HAS_DDCTD `i_axi_AXI_M12_SHARED_R_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M12_SHARED_B_HAS_DDCTD
  `define AXI_M12_SHARED_B_HAS_DDCTD `i_axi_AXI_M12_SHARED_B_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M13_SHARED_R_HAS_DDCTD
  `define AXI_M13_SHARED_R_HAS_DDCTD `i_axi_AXI_M13_SHARED_R_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M13_SHARED_B_HAS_DDCTD
  `define AXI_M13_SHARED_B_HAS_DDCTD `i_axi_AXI_M13_SHARED_B_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M14_SHARED_R_HAS_DDCTD
  `define AXI_M14_SHARED_R_HAS_DDCTD `i_axi_AXI_M14_SHARED_R_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M14_SHARED_B_HAS_DDCTD
  `define AXI_M14_SHARED_B_HAS_DDCTD `i_axi_AXI_M14_SHARED_B_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M15_SHARED_R_HAS_DDCTD
  `define AXI_M15_SHARED_R_HAS_DDCTD `i_axi_AXI_M15_SHARED_R_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_M15_SHARED_B_HAS_DDCTD
  `define AXI_M15_SHARED_B_HAS_DDCTD `i_axi_AXI_M15_SHARED_B_HAS_DDCTD
`endif 

`ifdef i_axi_AXI_PRIORITY_M1
  `define AXI_PRIORITY_M1 `i_axi_AXI_PRIORITY_M1
`endif 

`ifdef i_axi_AXI_PRIORITY_M2
  `define AXI_PRIORITY_M2 `i_axi_AXI_PRIORITY_M2
`endif 

`ifdef i_axi_AXI_PRIORITY_M3
  `define AXI_PRIORITY_M3 `i_axi_AXI_PRIORITY_M3
`endif 

`ifdef i_axi_AXI_PRIORITY_M4
  `define AXI_PRIORITY_M4 `i_axi_AXI_PRIORITY_M4
`endif 

`ifdef i_axi_AXI_PRIORITY_M5
  `define AXI_PRIORITY_M5 `i_axi_AXI_PRIORITY_M5
`endif 

`ifdef i_axi_AXI_PRIORITY_M6
  `define AXI_PRIORITY_M6 `i_axi_AXI_PRIORITY_M6
`endif 

`ifdef i_axi_AXI_PRIORITY_M7
  `define AXI_PRIORITY_M7 `i_axi_AXI_PRIORITY_M7
`endif 

`ifdef i_axi_AXI_PRIORITY_M8
  `define AXI_PRIORITY_M8 `i_axi_AXI_PRIORITY_M8
`endif 

`ifdef i_axi_AXI_PRIORITY_M9
  `define AXI_PRIORITY_M9 `i_axi_AXI_PRIORITY_M9
`endif 

`ifdef i_axi_AXI_PRIORITY_M10
  `define AXI_PRIORITY_M10 `i_axi_AXI_PRIORITY_M10
`endif 

`ifdef i_axi_AXI_PRIORITY_M11
  `define AXI_PRIORITY_M11 `i_axi_AXI_PRIORITY_M11
`endif 

`ifdef i_axi_AXI_PRIORITY_M12
  `define AXI_PRIORITY_M12 `i_axi_AXI_PRIORITY_M12
`endif 

`ifdef i_axi_AXI_PRIORITY_M13
  `define AXI_PRIORITY_M13 `i_axi_AXI_PRIORITY_M13
`endif 

`ifdef i_axi_AXI_PRIORITY_M14
  `define AXI_PRIORITY_M14 `i_axi_AXI_PRIORITY_M14
`endif 

`ifdef i_axi_AXI_PRIORITY_M15
  `define AXI_PRIORITY_M15 `i_axi_AXI_PRIORITY_M15
`endif 

`ifdef i_axi_AXI_PRIORITY_M16
  `define AXI_PRIORITY_M16 `i_axi_AXI_PRIORITY_M16
`endif 

`ifdef i_axi_AXI_PRIORITY_S1
  `define AXI_PRIORITY_S1 `i_axi_AXI_PRIORITY_S1
`endif 

`ifdef i_axi_AXI_PRIORITY_S2
  `define AXI_PRIORITY_S2 `i_axi_AXI_PRIORITY_S2
`endif 

`ifdef i_axi_AXI_PRIORITY_S3
  `define AXI_PRIORITY_S3 `i_axi_AXI_PRIORITY_S3
`endif 

`ifdef i_axi_AXI_PRIORITY_S4
  `define AXI_PRIORITY_S4 `i_axi_AXI_PRIORITY_S4
`endif 

`ifdef i_axi_AXI_PRIORITY_S5
  `define AXI_PRIORITY_S5 `i_axi_AXI_PRIORITY_S5
`endif 

`ifdef i_axi_AXI_PRIORITY_S6
  `define AXI_PRIORITY_S6 `i_axi_AXI_PRIORITY_S6
`endif 

`ifdef i_axi_AXI_PRIORITY_S7
  `define AXI_PRIORITY_S7 `i_axi_AXI_PRIORITY_S7
`endif 

`ifdef i_axi_AXI_PRIORITY_S8
  `define AXI_PRIORITY_S8 `i_axi_AXI_PRIORITY_S8
`endif 

`ifdef i_axi_AXI_PRIORITY_S9
  `define AXI_PRIORITY_S9 `i_axi_AXI_PRIORITY_S9
`endif 

`ifdef i_axi_AXI_PRIORITY_S10
  `define AXI_PRIORITY_S10 `i_axi_AXI_PRIORITY_S10
`endif 

`ifdef i_axi_AXI_PRIORITY_S11
  `define AXI_PRIORITY_S11 `i_axi_AXI_PRIORITY_S11
`endif 

`ifdef i_axi_AXI_PRIORITY_S12
  `define AXI_PRIORITY_S12 `i_axi_AXI_PRIORITY_S12
`endif 

`ifdef i_axi_AXI_PRIORITY_S13
  `define AXI_PRIORITY_S13 `i_axi_AXI_PRIORITY_S13
`endif 

`ifdef i_axi_AXI_PRIORITY_S14
  `define AXI_PRIORITY_S14 `i_axi_AXI_PRIORITY_S14
`endif 

`ifdef i_axi_AXI_PRIORITY_S15
  `define AXI_PRIORITY_S15 `i_axi_AXI_PRIORITY_S15
`endif 

`ifdef i_axi_AXI_PRIORITY_S16
  `define AXI_PRIORITY_S16 `i_axi_AXI_PRIORITY_S16
`endif 

`ifdef i_axi_AXI_PRIORITY_S0
  `define AXI_PRIORITY_S0 `i_axi_AXI_PRIORITY_S0
`endif 

`ifdef i_axi_AXI_HAS_EXT_PRIORITY
  `define AXI_HAS_EXT_PRIORITY `i_axi_AXI_HAS_EXT_PRIORITY
`endif 

`ifdef i_axi_AXI_SHARED_LAYER_MASTER_PRIORITY_EN_VAL
  `define AXI_SHARED_LAYER_MASTER_PRIORITY_EN_VAL `i_axi_AXI_SHARED_LAYER_MASTER_PRIORITY_EN_VAL
`endif 

`ifdef i_axi_AXI_SHARED_LAYER_MASTER_PRIORITY_EN
  `define AXI_SHARED_LAYER_MASTER_PRIORITY_EN `i_axi_AXI_SHARED_LAYER_MASTER_PRIORITY_EN
`endif 

`ifdef i_axi_AXI_SHARED_LAYER_MASTER_PRIORITY
  `define AXI_SHARED_LAYER_MASTER_PRIORITY `i_axi_AXI_SHARED_LAYER_MASTER_PRIORITY
`endif 

`ifdef i_axi_AXI_SHARED_LAYER_SLAVE_PRIORITY_EN_VAL
  `define AXI_SHARED_LAYER_SLAVE_PRIORITY_EN_VAL `i_axi_AXI_SHARED_LAYER_SLAVE_PRIORITY_EN_VAL
`endif 

`ifdef i_axi_AXI_SHARED_LAYER_SLAVE_PRIORITY_EN
  `define AXI_SHARED_LAYER_SLAVE_PRIORITY_EN `i_axi_AXI_SHARED_LAYER_SLAVE_PRIORITY_EN
`endif 

`ifdef i_axi_AXI_SHARED_LAYER_SLAVE_PRIORITY
  `define AXI_SHARED_LAYER_SLAVE_PRIORITY `i_axi_AXI_SHARED_LAYER_SLAVE_PRIORITY
`endif 

`ifdef i_axi_AXI_AR_ARB_TYPE_S0
  `define AXI_AR_ARB_TYPE_S0 `i_axi_AXI_AR_ARB_TYPE_S0
`endif 

`ifdef i_axi_AXI_AW_ARB_TYPE_S0
  `define AXI_AW_ARB_TYPE_S0 `i_axi_AXI_AW_ARB_TYPE_S0
`endif 

`ifdef i_axi_AXI_AR_ARB_TYPE_S1
  `define AXI_AR_ARB_TYPE_S1 `i_axi_AXI_AR_ARB_TYPE_S1
`endif 

`ifdef i_axi_AXI_AW_ARB_TYPE_S1
  `define AXI_AW_ARB_TYPE_S1 `i_axi_AXI_AW_ARB_TYPE_S1
`endif 

`ifdef i_axi_AXI_AR_ARB_TYPE_S2
  `define AXI_AR_ARB_TYPE_S2 `i_axi_AXI_AR_ARB_TYPE_S2
`endif 

`ifdef i_axi_AXI_AW_ARB_TYPE_S2
  `define AXI_AW_ARB_TYPE_S2 `i_axi_AXI_AW_ARB_TYPE_S2
`endif 

`ifdef i_axi_AXI_AR_ARB_TYPE_S3
  `define AXI_AR_ARB_TYPE_S3 `i_axi_AXI_AR_ARB_TYPE_S3
`endif 

`ifdef i_axi_AXI_AW_ARB_TYPE_S3
  `define AXI_AW_ARB_TYPE_S3 `i_axi_AXI_AW_ARB_TYPE_S3
`endif 

`ifdef i_axi_AXI_AR_ARB_TYPE_S4
  `define AXI_AR_ARB_TYPE_S4 `i_axi_AXI_AR_ARB_TYPE_S4
`endif 

`ifdef i_axi_AXI_AW_ARB_TYPE_S4
  `define AXI_AW_ARB_TYPE_S4 `i_axi_AXI_AW_ARB_TYPE_S4
`endif 

`ifdef i_axi_AXI_AR_ARB_TYPE_S5
  `define AXI_AR_ARB_TYPE_S5 `i_axi_AXI_AR_ARB_TYPE_S5
`endif 

`ifdef i_axi_AXI_AW_ARB_TYPE_S5
  `define AXI_AW_ARB_TYPE_S5 `i_axi_AXI_AW_ARB_TYPE_S5
`endif 

`ifdef i_axi_AXI_AR_ARB_TYPE_S6
  `define AXI_AR_ARB_TYPE_S6 `i_axi_AXI_AR_ARB_TYPE_S6
`endif 

`ifdef i_axi_AXI_AW_ARB_TYPE_S6
  `define AXI_AW_ARB_TYPE_S6 `i_axi_AXI_AW_ARB_TYPE_S6
`endif 

`ifdef i_axi_AXI_AR_ARB_TYPE_S7
  `define AXI_AR_ARB_TYPE_S7 `i_axi_AXI_AR_ARB_TYPE_S7
`endif 

`ifdef i_axi_AXI_AW_ARB_TYPE_S7
  `define AXI_AW_ARB_TYPE_S7 `i_axi_AXI_AW_ARB_TYPE_S7
`endif 

`ifdef i_axi_AXI_AR_ARB_TYPE_S8
  `define AXI_AR_ARB_TYPE_S8 `i_axi_AXI_AR_ARB_TYPE_S8
`endif 

`ifdef i_axi_AXI_AW_ARB_TYPE_S8
  `define AXI_AW_ARB_TYPE_S8 `i_axi_AXI_AW_ARB_TYPE_S8
`endif 

`ifdef i_axi_AXI_AR_ARB_TYPE_S9
  `define AXI_AR_ARB_TYPE_S9 `i_axi_AXI_AR_ARB_TYPE_S9
`endif 

`ifdef i_axi_AXI_AW_ARB_TYPE_S9
  `define AXI_AW_ARB_TYPE_S9 `i_axi_AXI_AW_ARB_TYPE_S9
`endif 

`ifdef i_axi_AXI_AR_ARB_TYPE_S10
  `define AXI_AR_ARB_TYPE_S10 `i_axi_AXI_AR_ARB_TYPE_S10
`endif 

`ifdef i_axi_AXI_AW_ARB_TYPE_S10
  `define AXI_AW_ARB_TYPE_S10 `i_axi_AXI_AW_ARB_TYPE_S10
`endif 

`ifdef i_axi_AXI_AR_ARB_TYPE_S11
  `define AXI_AR_ARB_TYPE_S11 `i_axi_AXI_AR_ARB_TYPE_S11
`endif 

`ifdef i_axi_AXI_AW_ARB_TYPE_S11
  `define AXI_AW_ARB_TYPE_S11 `i_axi_AXI_AW_ARB_TYPE_S11
`endif 

`ifdef i_axi_AXI_AR_ARB_TYPE_S12
  `define AXI_AR_ARB_TYPE_S12 `i_axi_AXI_AR_ARB_TYPE_S12
`endif 

`ifdef i_axi_AXI_AW_ARB_TYPE_S12
  `define AXI_AW_ARB_TYPE_S12 `i_axi_AXI_AW_ARB_TYPE_S12
`endif 

`ifdef i_axi_AXI_AR_ARB_TYPE_S13
  `define AXI_AR_ARB_TYPE_S13 `i_axi_AXI_AR_ARB_TYPE_S13
`endif 

`ifdef i_axi_AXI_AW_ARB_TYPE_S13
  `define AXI_AW_ARB_TYPE_S13 `i_axi_AXI_AW_ARB_TYPE_S13
`endif 

`ifdef i_axi_AXI_AR_ARB_TYPE_S14
  `define AXI_AR_ARB_TYPE_S14 `i_axi_AXI_AR_ARB_TYPE_S14
`endif 

`ifdef i_axi_AXI_AW_ARB_TYPE_S14
  `define AXI_AW_ARB_TYPE_S14 `i_axi_AXI_AW_ARB_TYPE_S14
`endif 

`ifdef i_axi_AXI_AR_ARB_TYPE_S15
  `define AXI_AR_ARB_TYPE_S15 `i_axi_AXI_AR_ARB_TYPE_S15
`endif 

`ifdef i_axi_AXI_AW_ARB_TYPE_S15
  `define AXI_AW_ARB_TYPE_S15 `i_axi_AXI_AW_ARB_TYPE_S15
`endif 

`ifdef i_axi_AXI_AR_ARB_TYPE_S16
  `define AXI_AR_ARB_TYPE_S16 `i_axi_AXI_AR_ARB_TYPE_S16
`endif 

`ifdef i_axi_AXI_AW_ARB_TYPE_S16
  `define AXI_AW_ARB_TYPE_S16 `i_axi_AXI_AW_ARB_TYPE_S16
`endif 

`ifdef i_axi_AXI_W_ARB_TYPE_S0
  `define AXI_W_ARB_TYPE_S0 `i_axi_AXI_W_ARB_TYPE_S0
`endif 

`ifdef i_axi_AXI_W_ARB_TYPE_S1
  `define AXI_W_ARB_TYPE_S1 `i_axi_AXI_W_ARB_TYPE_S1
`endif 

`ifdef i_axi_AXI_W_ARB_TYPE_S2
  `define AXI_W_ARB_TYPE_S2 `i_axi_AXI_W_ARB_TYPE_S2
`endif 

`ifdef i_axi_AXI_W_ARB_TYPE_S3
  `define AXI_W_ARB_TYPE_S3 `i_axi_AXI_W_ARB_TYPE_S3
`endif 

`ifdef i_axi_AXI_W_ARB_TYPE_S4
  `define AXI_W_ARB_TYPE_S4 `i_axi_AXI_W_ARB_TYPE_S4
`endif 

`ifdef i_axi_AXI_W_ARB_TYPE_S5
  `define AXI_W_ARB_TYPE_S5 `i_axi_AXI_W_ARB_TYPE_S5
`endif 

`ifdef i_axi_AXI_W_ARB_TYPE_S6
  `define AXI_W_ARB_TYPE_S6 `i_axi_AXI_W_ARB_TYPE_S6
`endif 

`ifdef i_axi_AXI_W_ARB_TYPE_S7
  `define AXI_W_ARB_TYPE_S7 `i_axi_AXI_W_ARB_TYPE_S7
`endif 

`ifdef i_axi_AXI_W_ARB_TYPE_S8
  `define AXI_W_ARB_TYPE_S8 `i_axi_AXI_W_ARB_TYPE_S8
`endif 

`ifdef i_axi_AXI_W_ARB_TYPE_S9
  `define AXI_W_ARB_TYPE_S9 `i_axi_AXI_W_ARB_TYPE_S9
`endif 

`ifdef i_axi_AXI_W_ARB_TYPE_S10
  `define AXI_W_ARB_TYPE_S10 `i_axi_AXI_W_ARB_TYPE_S10
`endif 

`ifdef i_axi_AXI_W_ARB_TYPE_S11
  `define AXI_W_ARB_TYPE_S11 `i_axi_AXI_W_ARB_TYPE_S11
`endif 

`ifdef i_axi_AXI_W_ARB_TYPE_S12
  `define AXI_W_ARB_TYPE_S12 `i_axi_AXI_W_ARB_TYPE_S12
`endif 

`ifdef i_axi_AXI_W_ARB_TYPE_S13
  `define AXI_W_ARB_TYPE_S13 `i_axi_AXI_W_ARB_TYPE_S13
`endif 

`ifdef i_axi_AXI_W_ARB_TYPE_S14
  `define AXI_W_ARB_TYPE_S14 `i_axi_AXI_W_ARB_TYPE_S14
`endif 

`ifdef i_axi_AXI_W_ARB_TYPE_S15
  `define AXI_W_ARB_TYPE_S15 `i_axi_AXI_W_ARB_TYPE_S15
`endif 

`ifdef i_axi_AXI_W_ARB_TYPE_S16
  `define AXI_W_ARB_TYPE_S16 `i_axi_AXI_W_ARB_TYPE_S16
`endif 

`ifdef i_axi_AXI_R_ARB_TYPE_M1
  `define AXI_R_ARB_TYPE_M1 `i_axi_AXI_R_ARB_TYPE_M1
`endif 

`ifdef i_axi_AXI_B_ARB_TYPE_M1
  `define AXI_B_ARB_TYPE_M1 `i_axi_AXI_B_ARB_TYPE_M1
`endif 

`ifdef i_axi_AXI_R_ARB_TYPE_M2
  `define AXI_R_ARB_TYPE_M2 `i_axi_AXI_R_ARB_TYPE_M2
`endif 

`ifdef i_axi_AXI_B_ARB_TYPE_M2
  `define AXI_B_ARB_TYPE_M2 `i_axi_AXI_B_ARB_TYPE_M2
`endif 

`ifdef i_axi_AXI_R_ARB_TYPE_M3
  `define AXI_R_ARB_TYPE_M3 `i_axi_AXI_R_ARB_TYPE_M3
`endif 

`ifdef i_axi_AXI_B_ARB_TYPE_M3
  `define AXI_B_ARB_TYPE_M3 `i_axi_AXI_B_ARB_TYPE_M3
`endif 

`ifdef i_axi_AXI_R_ARB_TYPE_M4
  `define AXI_R_ARB_TYPE_M4 `i_axi_AXI_R_ARB_TYPE_M4
`endif 

`ifdef i_axi_AXI_B_ARB_TYPE_M4
  `define AXI_B_ARB_TYPE_M4 `i_axi_AXI_B_ARB_TYPE_M4
`endif 

`ifdef i_axi_AXI_R_ARB_TYPE_M5
  `define AXI_R_ARB_TYPE_M5 `i_axi_AXI_R_ARB_TYPE_M5
`endif 

`ifdef i_axi_AXI_B_ARB_TYPE_M5
  `define AXI_B_ARB_TYPE_M5 `i_axi_AXI_B_ARB_TYPE_M5
`endif 

`ifdef i_axi_AXI_R_ARB_TYPE_M6
  `define AXI_R_ARB_TYPE_M6 `i_axi_AXI_R_ARB_TYPE_M6
`endif 

`ifdef i_axi_AXI_B_ARB_TYPE_M6
  `define AXI_B_ARB_TYPE_M6 `i_axi_AXI_B_ARB_TYPE_M6
`endif 

`ifdef i_axi_AXI_R_ARB_TYPE_M7
  `define AXI_R_ARB_TYPE_M7 `i_axi_AXI_R_ARB_TYPE_M7
`endif 

`ifdef i_axi_AXI_B_ARB_TYPE_M7
  `define AXI_B_ARB_TYPE_M7 `i_axi_AXI_B_ARB_TYPE_M7
`endif 

`ifdef i_axi_AXI_R_ARB_TYPE_M8
  `define AXI_R_ARB_TYPE_M8 `i_axi_AXI_R_ARB_TYPE_M8
`endif 

`ifdef i_axi_AXI_B_ARB_TYPE_M8
  `define AXI_B_ARB_TYPE_M8 `i_axi_AXI_B_ARB_TYPE_M8
`endif 

`ifdef i_axi_AXI_R_ARB_TYPE_M9
  `define AXI_R_ARB_TYPE_M9 `i_axi_AXI_R_ARB_TYPE_M9
`endif 

`ifdef i_axi_AXI_B_ARB_TYPE_M9
  `define AXI_B_ARB_TYPE_M9 `i_axi_AXI_B_ARB_TYPE_M9
`endif 

`ifdef i_axi_AXI_R_ARB_TYPE_M10
  `define AXI_R_ARB_TYPE_M10 `i_axi_AXI_R_ARB_TYPE_M10
`endif 

`ifdef i_axi_AXI_B_ARB_TYPE_M10
  `define AXI_B_ARB_TYPE_M10 `i_axi_AXI_B_ARB_TYPE_M10
`endif 

`ifdef i_axi_AXI_R_ARB_TYPE_M11
  `define AXI_R_ARB_TYPE_M11 `i_axi_AXI_R_ARB_TYPE_M11
`endif 

`ifdef i_axi_AXI_B_ARB_TYPE_M11
  `define AXI_B_ARB_TYPE_M11 `i_axi_AXI_B_ARB_TYPE_M11
`endif 

`ifdef i_axi_AXI_R_ARB_TYPE_M12
  `define AXI_R_ARB_TYPE_M12 `i_axi_AXI_R_ARB_TYPE_M12
`endif 

`ifdef i_axi_AXI_B_ARB_TYPE_M12
  `define AXI_B_ARB_TYPE_M12 `i_axi_AXI_B_ARB_TYPE_M12
`endif 

`ifdef i_axi_AXI_R_ARB_TYPE_M13
  `define AXI_R_ARB_TYPE_M13 `i_axi_AXI_R_ARB_TYPE_M13
`endif 

`ifdef i_axi_AXI_B_ARB_TYPE_M13
  `define AXI_B_ARB_TYPE_M13 `i_axi_AXI_B_ARB_TYPE_M13
`endif 

`ifdef i_axi_AXI_R_ARB_TYPE_M14
  `define AXI_R_ARB_TYPE_M14 `i_axi_AXI_R_ARB_TYPE_M14
`endif 

`ifdef i_axi_AXI_B_ARB_TYPE_M14
  `define AXI_B_ARB_TYPE_M14 `i_axi_AXI_B_ARB_TYPE_M14
`endif 

`ifdef i_axi_AXI_R_ARB_TYPE_M15
  `define AXI_R_ARB_TYPE_M15 `i_axi_AXI_R_ARB_TYPE_M15
`endif 

`ifdef i_axi_AXI_B_ARB_TYPE_M15
  `define AXI_B_ARB_TYPE_M15 `i_axi_AXI_B_ARB_TYPE_M15
`endif 

`ifdef i_axi_AXI_R_ARB_TYPE_M16
  `define AXI_R_ARB_TYPE_M16 `i_axi_AXI_R_ARB_TYPE_M16
`endif 

`ifdef i_axi_AXI_B_ARB_TYPE_M16
  `define AXI_B_ARB_TYPE_M16 `i_axi_AXI_B_ARB_TYPE_M16
`endif 

`ifdef i_axi_AXI_AR_SHARED_ARB_TYPE
  `define AXI_AR_SHARED_ARB_TYPE `i_axi_AXI_AR_SHARED_ARB_TYPE
`endif 

`ifdef i_axi_AXI_AW_SHARED_ARB_TYPE
  `define AXI_AW_SHARED_ARB_TYPE `i_axi_AXI_AW_SHARED_ARB_TYPE
`endif 

`ifdef i_axi_AXI_W_SHARED_ARB_TYPE
  `define AXI_W_SHARED_ARB_TYPE `i_axi_AXI_W_SHARED_ARB_TYPE
`endif 

`ifdef i_axi_AXI_R_SHARED_ARB_TYPE
  `define AXI_R_SHARED_ARB_TYPE `i_axi_AXI_R_SHARED_ARB_TYPE
`endif 

`ifdef i_axi_AXI_B_SHARED_ARB_TYPE
  `define AXI_B_SHARED_ARB_TYPE `i_axi_AXI_B_SHARED_ARB_TYPE
`endif 

`ifdef i_axi_AXI_USER_ARB_REMOVAL
  `define AXI_USER_ARB_REMOVAL `i_axi_AXI_USER_ARB_REMOVAL
`endif 

`ifdef i_axi_AXI_NUM_RN_S1
  `define AXI_NUM_RN_S1 `i_axi_AXI_NUM_RN_S1
`endif 

`ifdef i_axi_AXI_NUM_RN_S2
  `define AXI_NUM_RN_S2 `i_axi_AXI_NUM_RN_S2
`endif 

`ifdef i_axi_AXI_NUM_RN_S3
  `define AXI_NUM_RN_S3 `i_axi_AXI_NUM_RN_S3
`endif 

`ifdef i_axi_AXI_NUM_RN_S4
  `define AXI_NUM_RN_S4 `i_axi_AXI_NUM_RN_S4
`endif 

`ifdef i_axi_AXI_NUM_RN_S5
  `define AXI_NUM_RN_S5 `i_axi_AXI_NUM_RN_S5
`endif 

`ifdef i_axi_AXI_NUM_RN_S6
  `define AXI_NUM_RN_S6 `i_axi_AXI_NUM_RN_S6
`endif 

`ifdef i_axi_AXI_NUM_RN_S7
  `define AXI_NUM_RN_S7 `i_axi_AXI_NUM_RN_S7
`endif 

`ifdef i_axi_AXI_NUM_RN_S8
  `define AXI_NUM_RN_S8 `i_axi_AXI_NUM_RN_S8
`endif 

`ifdef i_axi_AXI_NUM_RN_S9
  `define AXI_NUM_RN_S9 `i_axi_AXI_NUM_RN_S9
`endif 

`ifdef i_axi_AXI_NUM_RN_S10
  `define AXI_NUM_RN_S10 `i_axi_AXI_NUM_RN_S10
`endif 

`ifdef i_axi_AXI_NUM_RN_S11
  `define AXI_NUM_RN_S11 `i_axi_AXI_NUM_RN_S11
`endif 

`ifdef i_axi_AXI_NUM_RN_S12
  `define AXI_NUM_RN_S12 `i_axi_AXI_NUM_RN_S12
`endif 

`ifdef i_axi_AXI_NUM_RN_S13
  `define AXI_NUM_RN_S13 `i_axi_AXI_NUM_RN_S13
`endif 

`ifdef i_axi_AXI_NUM_RN_S14
  `define AXI_NUM_RN_S14 `i_axi_AXI_NUM_RN_S14
`endif 

`ifdef i_axi_AXI_NUM_RN_S15
  `define AXI_NUM_RN_S15 `i_axi_AXI_NUM_RN_S15
`endif 

`ifdef i_axi_AXI_NUM_RN_S16
  `define AXI_NUM_RN_S16 `i_axi_AXI_NUM_RN_S16
`endif 

`ifdef i_axi_AXI_R1_NSA_S1
  `define AXI_R1_NSA_S1 `i_axi_AXI_R1_NSA_S1
`endif 

`ifdef i_axi_AXI_R1_NEA_S1
  `define AXI_R1_NEA_S1 `i_axi_AXI_R1_NEA_S1
`endif 

`ifdef i_axi_AXI_R1_NSA_S2
  `define AXI_R1_NSA_S2 `i_axi_AXI_R1_NSA_S2
`endif 

`ifdef i_axi_AXI_R1_NEA_S2
  `define AXI_R1_NEA_S2 `i_axi_AXI_R1_NEA_S2
`endif 

`ifdef i_axi_AXI_R1_NSA_S3
  `define AXI_R1_NSA_S3 `i_axi_AXI_R1_NSA_S3
`endif 

`ifdef i_axi_AXI_R1_NEA_S3
  `define AXI_R1_NEA_S3 `i_axi_AXI_R1_NEA_S3
`endif 

`ifdef i_axi_AXI_R1_NSA_S4
  `define AXI_R1_NSA_S4 `i_axi_AXI_R1_NSA_S4
`endif 

`ifdef i_axi_AXI_R1_NEA_S4
  `define AXI_R1_NEA_S4 `i_axi_AXI_R1_NEA_S4
`endif 

`ifdef i_axi_AXI_R1_NSA_S5
  `define AXI_R1_NSA_S5 `i_axi_AXI_R1_NSA_S5
`endif 

`ifdef i_axi_AXI_R1_NEA_S5
  `define AXI_R1_NEA_S5 `i_axi_AXI_R1_NEA_S5
`endif 

`ifdef i_axi_AXI_R1_NSA_S6
  `define AXI_R1_NSA_S6 `i_axi_AXI_R1_NSA_S6
`endif 

`ifdef i_axi_AXI_R1_NEA_S6
  `define AXI_R1_NEA_S6 `i_axi_AXI_R1_NEA_S6
`endif 

`ifdef i_axi_AXI_R1_NSA_S7
  `define AXI_R1_NSA_S7 `i_axi_AXI_R1_NSA_S7
`endif 

`ifdef i_axi_AXI_R1_NEA_S7
  `define AXI_R1_NEA_S7 `i_axi_AXI_R1_NEA_S7
`endif 

`ifdef i_axi_AXI_R1_NSA_S8
  `define AXI_R1_NSA_S8 `i_axi_AXI_R1_NSA_S8
`endif 

`ifdef i_axi_AXI_R1_NEA_S8
  `define AXI_R1_NEA_S8 `i_axi_AXI_R1_NEA_S8
`endif 

`ifdef i_axi_AXI_R1_NSA_S9
  `define AXI_R1_NSA_S9 `i_axi_AXI_R1_NSA_S9
`endif 

`ifdef i_axi_AXI_R1_NEA_S9
  `define AXI_R1_NEA_S9 `i_axi_AXI_R1_NEA_S9
`endif 

`ifdef i_axi_AXI_R1_NSA_S10
  `define AXI_R1_NSA_S10 `i_axi_AXI_R1_NSA_S10
`endif 

`ifdef i_axi_AXI_R1_NEA_S10
  `define AXI_R1_NEA_S10 `i_axi_AXI_R1_NEA_S10
`endif 

`ifdef i_axi_AXI_R1_NSA_S11
  `define AXI_R1_NSA_S11 `i_axi_AXI_R1_NSA_S11
`endif 

`ifdef i_axi_AXI_R1_NEA_S11
  `define AXI_R1_NEA_S11 `i_axi_AXI_R1_NEA_S11
`endif 

`ifdef i_axi_AXI_R1_NSA_S12
  `define AXI_R1_NSA_S12 `i_axi_AXI_R1_NSA_S12
`endif 

`ifdef i_axi_AXI_R1_NEA_S12
  `define AXI_R1_NEA_S12 `i_axi_AXI_R1_NEA_S12
`endif 

`ifdef i_axi_AXI_R1_NSA_S13
  `define AXI_R1_NSA_S13 `i_axi_AXI_R1_NSA_S13
`endif 

`ifdef i_axi_AXI_R1_NEA_S13
  `define AXI_R1_NEA_S13 `i_axi_AXI_R1_NEA_S13
`endif 

`ifdef i_axi_AXI_R1_NSA_S14
  `define AXI_R1_NSA_S14 `i_axi_AXI_R1_NSA_S14
`endif 

`ifdef i_axi_AXI_R1_NEA_S14
  `define AXI_R1_NEA_S14 `i_axi_AXI_R1_NEA_S14
`endif 

`ifdef i_axi_AXI_R1_NSA_S15
  `define AXI_R1_NSA_S15 `i_axi_AXI_R1_NSA_S15
`endif 

`ifdef i_axi_AXI_R1_NEA_S15
  `define AXI_R1_NEA_S15 `i_axi_AXI_R1_NEA_S15
`endif 

`ifdef i_axi_AXI_R1_NSA_S16
  `define AXI_R1_NSA_S16 `i_axi_AXI_R1_NSA_S16
`endif 

`ifdef i_axi_AXI_R1_NEA_S16
  `define AXI_R1_NEA_S16 `i_axi_AXI_R1_NEA_S16
`endif 

`ifdef i_axi_AXI_R2_NSA_S1
  `define AXI_R2_NSA_S1 `i_axi_AXI_R2_NSA_S1
`endif 

`ifdef i_axi_AXI_R2_NEA_S1
  `define AXI_R2_NEA_S1 `i_axi_AXI_R2_NEA_S1
`endif 

`ifdef i_axi_AXI_R2_NSA_S2
  `define AXI_R2_NSA_S2 `i_axi_AXI_R2_NSA_S2
`endif 

`ifdef i_axi_AXI_R2_NEA_S2
  `define AXI_R2_NEA_S2 `i_axi_AXI_R2_NEA_S2
`endif 

`ifdef i_axi_AXI_R2_NSA_S3
  `define AXI_R2_NSA_S3 `i_axi_AXI_R2_NSA_S3
`endif 

`ifdef i_axi_AXI_R2_NEA_S3
  `define AXI_R2_NEA_S3 `i_axi_AXI_R2_NEA_S3
`endif 

`ifdef i_axi_AXI_R2_NSA_S4
  `define AXI_R2_NSA_S4 `i_axi_AXI_R2_NSA_S4
`endif 

`ifdef i_axi_AXI_R2_NEA_S4
  `define AXI_R2_NEA_S4 `i_axi_AXI_R2_NEA_S4
`endif 

`ifdef i_axi_AXI_R2_NSA_S5
  `define AXI_R2_NSA_S5 `i_axi_AXI_R2_NSA_S5
`endif 

`ifdef i_axi_AXI_R2_NEA_S5
  `define AXI_R2_NEA_S5 `i_axi_AXI_R2_NEA_S5
`endif 

`ifdef i_axi_AXI_R2_NSA_S6
  `define AXI_R2_NSA_S6 `i_axi_AXI_R2_NSA_S6
`endif 

`ifdef i_axi_AXI_R2_NEA_S6
  `define AXI_R2_NEA_S6 `i_axi_AXI_R2_NEA_S6
`endif 

`ifdef i_axi_AXI_R2_NSA_S7
  `define AXI_R2_NSA_S7 `i_axi_AXI_R2_NSA_S7
`endif 

`ifdef i_axi_AXI_R2_NEA_S7
  `define AXI_R2_NEA_S7 `i_axi_AXI_R2_NEA_S7
`endif 

`ifdef i_axi_AXI_R2_NSA_S8
  `define AXI_R2_NSA_S8 `i_axi_AXI_R2_NSA_S8
`endif 

`ifdef i_axi_AXI_R2_NEA_S8
  `define AXI_R2_NEA_S8 `i_axi_AXI_R2_NEA_S8
`endif 

`ifdef i_axi_AXI_R2_NSA_S9
  `define AXI_R2_NSA_S9 `i_axi_AXI_R2_NSA_S9
`endif 

`ifdef i_axi_AXI_R2_NEA_S9
  `define AXI_R2_NEA_S9 `i_axi_AXI_R2_NEA_S9
`endif 

`ifdef i_axi_AXI_R2_NSA_S10
  `define AXI_R2_NSA_S10 `i_axi_AXI_R2_NSA_S10
`endif 

`ifdef i_axi_AXI_R2_NEA_S10
  `define AXI_R2_NEA_S10 `i_axi_AXI_R2_NEA_S10
`endif 

`ifdef i_axi_AXI_R2_NSA_S11
  `define AXI_R2_NSA_S11 `i_axi_AXI_R2_NSA_S11
`endif 

`ifdef i_axi_AXI_R2_NEA_S11
  `define AXI_R2_NEA_S11 `i_axi_AXI_R2_NEA_S11
`endif 

`ifdef i_axi_AXI_R2_NSA_S12
  `define AXI_R2_NSA_S12 `i_axi_AXI_R2_NSA_S12
`endif 

`ifdef i_axi_AXI_R2_NEA_S12
  `define AXI_R2_NEA_S12 `i_axi_AXI_R2_NEA_S12
`endif 

`ifdef i_axi_AXI_R2_NSA_S13
  `define AXI_R2_NSA_S13 `i_axi_AXI_R2_NSA_S13
`endif 

`ifdef i_axi_AXI_R2_NEA_S13
  `define AXI_R2_NEA_S13 `i_axi_AXI_R2_NEA_S13
`endif 

`ifdef i_axi_AXI_R2_NSA_S14
  `define AXI_R2_NSA_S14 `i_axi_AXI_R2_NSA_S14
`endif 

`ifdef i_axi_AXI_R2_NEA_S14
  `define AXI_R2_NEA_S14 `i_axi_AXI_R2_NEA_S14
`endif 

`ifdef i_axi_AXI_R2_NSA_S15
  `define AXI_R2_NSA_S15 `i_axi_AXI_R2_NSA_S15
`endif 

`ifdef i_axi_AXI_R2_NEA_S15
  `define AXI_R2_NEA_S15 `i_axi_AXI_R2_NEA_S15
`endif 

`ifdef i_axi_AXI_R2_NSA_S16
  `define AXI_R2_NSA_S16 `i_axi_AXI_R2_NSA_S16
`endif 

`ifdef i_axi_AXI_R2_NEA_S16
  `define AXI_R2_NEA_S16 `i_axi_AXI_R2_NEA_S16
`endif 

`ifdef i_axi_AXI_R3_NSA_S1
  `define AXI_R3_NSA_S1 `i_axi_AXI_R3_NSA_S1
`endif 

`ifdef i_axi_AXI_R3_NEA_S1
  `define AXI_R3_NEA_S1 `i_axi_AXI_R3_NEA_S1
`endif 

`ifdef i_axi_AXI_R3_NSA_S2
  `define AXI_R3_NSA_S2 `i_axi_AXI_R3_NSA_S2
`endif 

`ifdef i_axi_AXI_R3_NEA_S2
  `define AXI_R3_NEA_S2 `i_axi_AXI_R3_NEA_S2
`endif 

`ifdef i_axi_AXI_R3_NSA_S3
  `define AXI_R3_NSA_S3 `i_axi_AXI_R3_NSA_S3
`endif 

`ifdef i_axi_AXI_R3_NEA_S3
  `define AXI_R3_NEA_S3 `i_axi_AXI_R3_NEA_S3
`endif 

`ifdef i_axi_AXI_R3_NSA_S4
  `define AXI_R3_NSA_S4 `i_axi_AXI_R3_NSA_S4
`endif 

`ifdef i_axi_AXI_R3_NEA_S4
  `define AXI_R3_NEA_S4 `i_axi_AXI_R3_NEA_S4
`endif 

`ifdef i_axi_AXI_R3_NSA_S5
  `define AXI_R3_NSA_S5 `i_axi_AXI_R3_NSA_S5
`endif 

`ifdef i_axi_AXI_R3_NEA_S5
  `define AXI_R3_NEA_S5 `i_axi_AXI_R3_NEA_S5
`endif 

`ifdef i_axi_AXI_R3_NSA_S6
  `define AXI_R3_NSA_S6 `i_axi_AXI_R3_NSA_S6
`endif 

`ifdef i_axi_AXI_R3_NEA_S6
  `define AXI_R3_NEA_S6 `i_axi_AXI_R3_NEA_S6
`endif 

`ifdef i_axi_AXI_R3_NSA_S7
  `define AXI_R3_NSA_S7 `i_axi_AXI_R3_NSA_S7
`endif 

`ifdef i_axi_AXI_R3_NEA_S7
  `define AXI_R3_NEA_S7 `i_axi_AXI_R3_NEA_S7
`endif 

`ifdef i_axi_AXI_R3_NSA_S8
  `define AXI_R3_NSA_S8 `i_axi_AXI_R3_NSA_S8
`endif 

`ifdef i_axi_AXI_R3_NEA_S8
  `define AXI_R3_NEA_S8 `i_axi_AXI_R3_NEA_S8
`endif 

`ifdef i_axi_AXI_R3_NSA_S9
  `define AXI_R3_NSA_S9 `i_axi_AXI_R3_NSA_S9
`endif 

`ifdef i_axi_AXI_R3_NEA_S9
  `define AXI_R3_NEA_S9 `i_axi_AXI_R3_NEA_S9
`endif 

`ifdef i_axi_AXI_R3_NSA_S10
  `define AXI_R3_NSA_S10 `i_axi_AXI_R3_NSA_S10
`endif 

`ifdef i_axi_AXI_R3_NEA_S10
  `define AXI_R3_NEA_S10 `i_axi_AXI_R3_NEA_S10
`endif 

`ifdef i_axi_AXI_R3_NSA_S11
  `define AXI_R3_NSA_S11 `i_axi_AXI_R3_NSA_S11
`endif 

`ifdef i_axi_AXI_R3_NEA_S11
  `define AXI_R3_NEA_S11 `i_axi_AXI_R3_NEA_S11
`endif 

`ifdef i_axi_AXI_R3_NSA_S12
  `define AXI_R3_NSA_S12 `i_axi_AXI_R3_NSA_S12
`endif 

`ifdef i_axi_AXI_R3_NEA_S12
  `define AXI_R3_NEA_S12 `i_axi_AXI_R3_NEA_S12
`endif 

`ifdef i_axi_AXI_R3_NSA_S13
  `define AXI_R3_NSA_S13 `i_axi_AXI_R3_NSA_S13
`endif 

`ifdef i_axi_AXI_R3_NEA_S13
  `define AXI_R3_NEA_S13 `i_axi_AXI_R3_NEA_S13
`endif 

`ifdef i_axi_AXI_R3_NSA_S14
  `define AXI_R3_NSA_S14 `i_axi_AXI_R3_NSA_S14
`endif 

`ifdef i_axi_AXI_R3_NEA_S14
  `define AXI_R3_NEA_S14 `i_axi_AXI_R3_NEA_S14
`endif 

`ifdef i_axi_AXI_R3_NSA_S15
  `define AXI_R3_NSA_S15 `i_axi_AXI_R3_NSA_S15
`endif 

`ifdef i_axi_AXI_R3_NEA_S15
  `define AXI_R3_NEA_S15 `i_axi_AXI_R3_NEA_S15
`endif 

`ifdef i_axi_AXI_R3_NSA_S16
  `define AXI_R3_NSA_S16 `i_axi_AXI_R3_NSA_S16
`endif 

`ifdef i_axi_AXI_R3_NEA_S16
  `define AXI_R3_NEA_S16 `i_axi_AXI_R3_NEA_S16
`endif 

`ifdef i_axi_AXI_R4_NSA_S1
  `define AXI_R4_NSA_S1 `i_axi_AXI_R4_NSA_S1
`endif 

`ifdef i_axi_AXI_R4_NEA_S1
  `define AXI_R4_NEA_S1 `i_axi_AXI_R4_NEA_S1
`endif 

`ifdef i_axi_AXI_R4_NSA_S2
  `define AXI_R4_NSA_S2 `i_axi_AXI_R4_NSA_S2
`endif 

`ifdef i_axi_AXI_R4_NEA_S2
  `define AXI_R4_NEA_S2 `i_axi_AXI_R4_NEA_S2
`endif 

`ifdef i_axi_AXI_R4_NSA_S3
  `define AXI_R4_NSA_S3 `i_axi_AXI_R4_NSA_S3
`endif 

`ifdef i_axi_AXI_R4_NEA_S3
  `define AXI_R4_NEA_S3 `i_axi_AXI_R4_NEA_S3
`endif 

`ifdef i_axi_AXI_R4_NSA_S4
  `define AXI_R4_NSA_S4 `i_axi_AXI_R4_NSA_S4
`endif 

`ifdef i_axi_AXI_R4_NEA_S4
  `define AXI_R4_NEA_S4 `i_axi_AXI_R4_NEA_S4
`endif 

`ifdef i_axi_AXI_R4_NSA_S5
  `define AXI_R4_NSA_S5 `i_axi_AXI_R4_NSA_S5
`endif 

`ifdef i_axi_AXI_R4_NEA_S5
  `define AXI_R4_NEA_S5 `i_axi_AXI_R4_NEA_S5
`endif 

`ifdef i_axi_AXI_R4_NSA_S6
  `define AXI_R4_NSA_S6 `i_axi_AXI_R4_NSA_S6
`endif 

`ifdef i_axi_AXI_R4_NEA_S6
  `define AXI_R4_NEA_S6 `i_axi_AXI_R4_NEA_S6
`endif 

`ifdef i_axi_AXI_R4_NSA_S7
  `define AXI_R4_NSA_S7 `i_axi_AXI_R4_NSA_S7
`endif 

`ifdef i_axi_AXI_R4_NEA_S7
  `define AXI_R4_NEA_S7 `i_axi_AXI_R4_NEA_S7
`endif 

`ifdef i_axi_AXI_R4_NSA_S8
  `define AXI_R4_NSA_S8 `i_axi_AXI_R4_NSA_S8
`endif 

`ifdef i_axi_AXI_R4_NEA_S8
  `define AXI_R4_NEA_S8 `i_axi_AXI_R4_NEA_S8
`endif 

`ifdef i_axi_AXI_R4_NSA_S9
  `define AXI_R4_NSA_S9 `i_axi_AXI_R4_NSA_S9
`endif 

`ifdef i_axi_AXI_R4_NEA_S9
  `define AXI_R4_NEA_S9 `i_axi_AXI_R4_NEA_S9
`endif 

`ifdef i_axi_AXI_R4_NSA_S10
  `define AXI_R4_NSA_S10 `i_axi_AXI_R4_NSA_S10
`endif 

`ifdef i_axi_AXI_R4_NEA_S10
  `define AXI_R4_NEA_S10 `i_axi_AXI_R4_NEA_S10
`endif 

`ifdef i_axi_AXI_R4_NSA_S11
  `define AXI_R4_NSA_S11 `i_axi_AXI_R4_NSA_S11
`endif 

`ifdef i_axi_AXI_R4_NEA_S11
  `define AXI_R4_NEA_S11 `i_axi_AXI_R4_NEA_S11
`endif 

`ifdef i_axi_AXI_R4_NSA_S12
  `define AXI_R4_NSA_S12 `i_axi_AXI_R4_NSA_S12
`endif 

`ifdef i_axi_AXI_R4_NEA_S12
  `define AXI_R4_NEA_S12 `i_axi_AXI_R4_NEA_S12
`endif 

`ifdef i_axi_AXI_R4_NSA_S13
  `define AXI_R4_NSA_S13 `i_axi_AXI_R4_NSA_S13
`endif 

`ifdef i_axi_AXI_R4_NEA_S13
  `define AXI_R4_NEA_S13 `i_axi_AXI_R4_NEA_S13
`endif 

`ifdef i_axi_AXI_R4_NSA_S14
  `define AXI_R4_NSA_S14 `i_axi_AXI_R4_NSA_S14
`endif 

`ifdef i_axi_AXI_R4_NEA_S14
  `define AXI_R4_NEA_S14 `i_axi_AXI_R4_NEA_S14
`endif 

`ifdef i_axi_AXI_R4_NSA_S15
  `define AXI_R4_NSA_S15 `i_axi_AXI_R4_NSA_S15
`endif 

`ifdef i_axi_AXI_R4_NEA_S15
  `define AXI_R4_NEA_S15 `i_axi_AXI_R4_NEA_S15
`endif 

`ifdef i_axi_AXI_R4_NSA_S16
  `define AXI_R4_NSA_S16 `i_axi_AXI_R4_NSA_S16
`endif 

`ifdef i_axi_AXI_R4_NEA_S16
  `define AXI_R4_NEA_S16 `i_axi_AXI_R4_NEA_S16
`endif 

`ifdef i_axi_AXI_R5_NSA_S1
  `define AXI_R5_NSA_S1 `i_axi_AXI_R5_NSA_S1
`endif 

`ifdef i_axi_AXI_R5_NEA_S1
  `define AXI_R5_NEA_S1 `i_axi_AXI_R5_NEA_S1
`endif 

`ifdef i_axi_AXI_R5_NSA_S2
  `define AXI_R5_NSA_S2 `i_axi_AXI_R5_NSA_S2
`endif 

`ifdef i_axi_AXI_R5_NEA_S2
  `define AXI_R5_NEA_S2 `i_axi_AXI_R5_NEA_S2
`endif 

`ifdef i_axi_AXI_R5_NSA_S3
  `define AXI_R5_NSA_S3 `i_axi_AXI_R5_NSA_S3
`endif 

`ifdef i_axi_AXI_R5_NEA_S3
  `define AXI_R5_NEA_S3 `i_axi_AXI_R5_NEA_S3
`endif 

`ifdef i_axi_AXI_R5_NSA_S4
  `define AXI_R5_NSA_S4 `i_axi_AXI_R5_NSA_S4
`endif 

`ifdef i_axi_AXI_R5_NEA_S4
  `define AXI_R5_NEA_S4 `i_axi_AXI_R5_NEA_S4
`endif 

`ifdef i_axi_AXI_R5_NSA_S5
  `define AXI_R5_NSA_S5 `i_axi_AXI_R5_NSA_S5
`endif 

`ifdef i_axi_AXI_R5_NEA_S5
  `define AXI_R5_NEA_S5 `i_axi_AXI_R5_NEA_S5
`endif 

`ifdef i_axi_AXI_R5_NSA_S6
  `define AXI_R5_NSA_S6 `i_axi_AXI_R5_NSA_S6
`endif 

`ifdef i_axi_AXI_R5_NEA_S6
  `define AXI_R5_NEA_S6 `i_axi_AXI_R5_NEA_S6
`endif 

`ifdef i_axi_AXI_R5_NSA_S7
  `define AXI_R5_NSA_S7 `i_axi_AXI_R5_NSA_S7
`endif 

`ifdef i_axi_AXI_R5_NEA_S7
  `define AXI_R5_NEA_S7 `i_axi_AXI_R5_NEA_S7
`endif 

`ifdef i_axi_AXI_R5_NSA_S8
  `define AXI_R5_NSA_S8 `i_axi_AXI_R5_NSA_S8
`endif 

`ifdef i_axi_AXI_R5_NEA_S8
  `define AXI_R5_NEA_S8 `i_axi_AXI_R5_NEA_S8
`endif 

`ifdef i_axi_AXI_R5_NSA_S9
  `define AXI_R5_NSA_S9 `i_axi_AXI_R5_NSA_S9
`endif 

`ifdef i_axi_AXI_R5_NEA_S9
  `define AXI_R5_NEA_S9 `i_axi_AXI_R5_NEA_S9
`endif 

`ifdef i_axi_AXI_R5_NSA_S10
  `define AXI_R5_NSA_S10 `i_axi_AXI_R5_NSA_S10
`endif 

`ifdef i_axi_AXI_R5_NEA_S10
  `define AXI_R5_NEA_S10 `i_axi_AXI_R5_NEA_S10
`endif 

`ifdef i_axi_AXI_R5_NSA_S11
  `define AXI_R5_NSA_S11 `i_axi_AXI_R5_NSA_S11
`endif 

`ifdef i_axi_AXI_R5_NEA_S11
  `define AXI_R5_NEA_S11 `i_axi_AXI_R5_NEA_S11
`endif 

`ifdef i_axi_AXI_R5_NSA_S12
  `define AXI_R5_NSA_S12 `i_axi_AXI_R5_NSA_S12
`endif 

`ifdef i_axi_AXI_R5_NEA_S12
  `define AXI_R5_NEA_S12 `i_axi_AXI_R5_NEA_S12
`endif 

`ifdef i_axi_AXI_R5_NSA_S13
  `define AXI_R5_NSA_S13 `i_axi_AXI_R5_NSA_S13
`endif 

`ifdef i_axi_AXI_R5_NEA_S13
  `define AXI_R5_NEA_S13 `i_axi_AXI_R5_NEA_S13
`endif 

`ifdef i_axi_AXI_R5_NSA_S14
  `define AXI_R5_NSA_S14 `i_axi_AXI_R5_NSA_S14
`endif 

`ifdef i_axi_AXI_R5_NEA_S14
  `define AXI_R5_NEA_S14 `i_axi_AXI_R5_NEA_S14
`endif 

`ifdef i_axi_AXI_R5_NSA_S15
  `define AXI_R5_NSA_S15 `i_axi_AXI_R5_NSA_S15
`endif 

`ifdef i_axi_AXI_R5_NEA_S15
  `define AXI_R5_NEA_S15 `i_axi_AXI_R5_NEA_S15
`endif 

`ifdef i_axi_AXI_R5_NSA_S16
  `define AXI_R5_NSA_S16 `i_axi_AXI_R5_NSA_S16
`endif 

`ifdef i_axi_AXI_R5_NEA_S16
  `define AXI_R5_NEA_S16 `i_axi_AXI_R5_NEA_S16
`endif 

`ifdef i_axi_AXI_R6_NSA_S1
  `define AXI_R6_NSA_S1 `i_axi_AXI_R6_NSA_S1
`endif 

`ifdef i_axi_AXI_R6_NEA_S1
  `define AXI_R6_NEA_S1 `i_axi_AXI_R6_NEA_S1
`endif 

`ifdef i_axi_AXI_R6_NSA_S2
  `define AXI_R6_NSA_S2 `i_axi_AXI_R6_NSA_S2
`endif 

`ifdef i_axi_AXI_R6_NEA_S2
  `define AXI_R6_NEA_S2 `i_axi_AXI_R6_NEA_S2
`endif 

`ifdef i_axi_AXI_R6_NSA_S3
  `define AXI_R6_NSA_S3 `i_axi_AXI_R6_NSA_S3
`endif 

`ifdef i_axi_AXI_R6_NEA_S3
  `define AXI_R6_NEA_S3 `i_axi_AXI_R6_NEA_S3
`endif 

`ifdef i_axi_AXI_R6_NSA_S4
  `define AXI_R6_NSA_S4 `i_axi_AXI_R6_NSA_S4
`endif 

`ifdef i_axi_AXI_R6_NEA_S4
  `define AXI_R6_NEA_S4 `i_axi_AXI_R6_NEA_S4
`endif 

`ifdef i_axi_AXI_R6_NSA_S5
  `define AXI_R6_NSA_S5 `i_axi_AXI_R6_NSA_S5
`endif 

`ifdef i_axi_AXI_R6_NEA_S5
  `define AXI_R6_NEA_S5 `i_axi_AXI_R6_NEA_S5
`endif 

`ifdef i_axi_AXI_R6_NSA_S6
  `define AXI_R6_NSA_S6 `i_axi_AXI_R6_NSA_S6
`endif 

`ifdef i_axi_AXI_R6_NEA_S6
  `define AXI_R6_NEA_S6 `i_axi_AXI_R6_NEA_S6
`endif 

`ifdef i_axi_AXI_R6_NSA_S7
  `define AXI_R6_NSA_S7 `i_axi_AXI_R6_NSA_S7
`endif 

`ifdef i_axi_AXI_R6_NEA_S7
  `define AXI_R6_NEA_S7 `i_axi_AXI_R6_NEA_S7
`endif 

`ifdef i_axi_AXI_R6_NSA_S8
  `define AXI_R6_NSA_S8 `i_axi_AXI_R6_NSA_S8
`endif 

`ifdef i_axi_AXI_R6_NEA_S8
  `define AXI_R6_NEA_S8 `i_axi_AXI_R6_NEA_S8
`endif 

`ifdef i_axi_AXI_R6_NSA_S9
  `define AXI_R6_NSA_S9 `i_axi_AXI_R6_NSA_S9
`endif 

`ifdef i_axi_AXI_R6_NEA_S9
  `define AXI_R6_NEA_S9 `i_axi_AXI_R6_NEA_S9
`endif 

`ifdef i_axi_AXI_R6_NSA_S10
  `define AXI_R6_NSA_S10 `i_axi_AXI_R6_NSA_S10
`endif 

`ifdef i_axi_AXI_R6_NEA_S10
  `define AXI_R6_NEA_S10 `i_axi_AXI_R6_NEA_S10
`endif 

`ifdef i_axi_AXI_R6_NSA_S11
  `define AXI_R6_NSA_S11 `i_axi_AXI_R6_NSA_S11
`endif 

`ifdef i_axi_AXI_R6_NEA_S11
  `define AXI_R6_NEA_S11 `i_axi_AXI_R6_NEA_S11
`endif 

`ifdef i_axi_AXI_R6_NSA_S12
  `define AXI_R6_NSA_S12 `i_axi_AXI_R6_NSA_S12
`endif 

`ifdef i_axi_AXI_R6_NEA_S12
  `define AXI_R6_NEA_S12 `i_axi_AXI_R6_NEA_S12
`endif 

`ifdef i_axi_AXI_R6_NSA_S13
  `define AXI_R6_NSA_S13 `i_axi_AXI_R6_NSA_S13
`endif 

`ifdef i_axi_AXI_R6_NEA_S13
  `define AXI_R6_NEA_S13 `i_axi_AXI_R6_NEA_S13
`endif 

`ifdef i_axi_AXI_R6_NSA_S14
  `define AXI_R6_NSA_S14 `i_axi_AXI_R6_NSA_S14
`endif 

`ifdef i_axi_AXI_R6_NEA_S14
  `define AXI_R6_NEA_S14 `i_axi_AXI_R6_NEA_S14
`endif 

`ifdef i_axi_AXI_R6_NSA_S15
  `define AXI_R6_NSA_S15 `i_axi_AXI_R6_NSA_S15
`endif 

`ifdef i_axi_AXI_R6_NEA_S15
  `define AXI_R6_NEA_S15 `i_axi_AXI_R6_NEA_S15
`endif 

`ifdef i_axi_AXI_R6_NSA_S16
  `define AXI_R6_NSA_S16 `i_axi_AXI_R6_NSA_S16
`endif 

`ifdef i_axi_AXI_R6_NEA_S16
  `define AXI_R6_NEA_S16 `i_axi_AXI_R6_NEA_S16
`endif 

`ifdef i_axi_AXI_R7_NSA_S1
  `define AXI_R7_NSA_S1 `i_axi_AXI_R7_NSA_S1
`endif 

`ifdef i_axi_AXI_R7_NEA_S1
  `define AXI_R7_NEA_S1 `i_axi_AXI_R7_NEA_S1
`endif 

`ifdef i_axi_AXI_R7_NSA_S2
  `define AXI_R7_NSA_S2 `i_axi_AXI_R7_NSA_S2
`endif 

`ifdef i_axi_AXI_R7_NEA_S2
  `define AXI_R7_NEA_S2 `i_axi_AXI_R7_NEA_S2
`endif 

`ifdef i_axi_AXI_R7_NSA_S3
  `define AXI_R7_NSA_S3 `i_axi_AXI_R7_NSA_S3
`endif 

`ifdef i_axi_AXI_R7_NEA_S3
  `define AXI_R7_NEA_S3 `i_axi_AXI_R7_NEA_S3
`endif 

`ifdef i_axi_AXI_R7_NSA_S4
  `define AXI_R7_NSA_S4 `i_axi_AXI_R7_NSA_S4
`endif 

`ifdef i_axi_AXI_R7_NEA_S4
  `define AXI_R7_NEA_S4 `i_axi_AXI_R7_NEA_S4
`endif 

`ifdef i_axi_AXI_R7_NSA_S5
  `define AXI_R7_NSA_S5 `i_axi_AXI_R7_NSA_S5
`endif 

`ifdef i_axi_AXI_R7_NEA_S5
  `define AXI_R7_NEA_S5 `i_axi_AXI_R7_NEA_S5
`endif 

`ifdef i_axi_AXI_R7_NSA_S6
  `define AXI_R7_NSA_S6 `i_axi_AXI_R7_NSA_S6
`endif 

`ifdef i_axi_AXI_R7_NEA_S6
  `define AXI_R7_NEA_S6 `i_axi_AXI_R7_NEA_S6
`endif 

`ifdef i_axi_AXI_R7_NSA_S7
  `define AXI_R7_NSA_S7 `i_axi_AXI_R7_NSA_S7
`endif 

`ifdef i_axi_AXI_R7_NEA_S7
  `define AXI_R7_NEA_S7 `i_axi_AXI_R7_NEA_S7
`endif 

`ifdef i_axi_AXI_R7_NSA_S8
  `define AXI_R7_NSA_S8 `i_axi_AXI_R7_NSA_S8
`endif 

`ifdef i_axi_AXI_R7_NEA_S8
  `define AXI_R7_NEA_S8 `i_axi_AXI_R7_NEA_S8
`endif 

`ifdef i_axi_AXI_R7_NSA_S9
  `define AXI_R7_NSA_S9 `i_axi_AXI_R7_NSA_S9
`endif 

`ifdef i_axi_AXI_R7_NEA_S9
  `define AXI_R7_NEA_S9 `i_axi_AXI_R7_NEA_S9
`endif 

`ifdef i_axi_AXI_R7_NSA_S10
  `define AXI_R7_NSA_S10 `i_axi_AXI_R7_NSA_S10
`endif 

`ifdef i_axi_AXI_R7_NEA_S10
  `define AXI_R7_NEA_S10 `i_axi_AXI_R7_NEA_S10
`endif 

`ifdef i_axi_AXI_R7_NSA_S11
  `define AXI_R7_NSA_S11 `i_axi_AXI_R7_NSA_S11
`endif 

`ifdef i_axi_AXI_R7_NEA_S11
  `define AXI_R7_NEA_S11 `i_axi_AXI_R7_NEA_S11
`endif 

`ifdef i_axi_AXI_R7_NSA_S12
  `define AXI_R7_NSA_S12 `i_axi_AXI_R7_NSA_S12
`endif 

`ifdef i_axi_AXI_R7_NEA_S12
  `define AXI_R7_NEA_S12 `i_axi_AXI_R7_NEA_S12
`endif 

`ifdef i_axi_AXI_R7_NSA_S13
  `define AXI_R7_NSA_S13 `i_axi_AXI_R7_NSA_S13
`endif 

`ifdef i_axi_AXI_R7_NEA_S13
  `define AXI_R7_NEA_S13 `i_axi_AXI_R7_NEA_S13
`endif 

`ifdef i_axi_AXI_R7_NSA_S14
  `define AXI_R7_NSA_S14 `i_axi_AXI_R7_NSA_S14
`endif 

`ifdef i_axi_AXI_R7_NEA_S14
  `define AXI_R7_NEA_S14 `i_axi_AXI_R7_NEA_S14
`endif 

`ifdef i_axi_AXI_R7_NSA_S15
  `define AXI_R7_NSA_S15 `i_axi_AXI_R7_NSA_S15
`endif 

`ifdef i_axi_AXI_R7_NEA_S15
  `define AXI_R7_NEA_S15 `i_axi_AXI_R7_NEA_S15
`endif 

`ifdef i_axi_AXI_R7_NSA_S16
  `define AXI_R7_NSA_S16 `i_axi_AXI_R7_NSA_S16
`endif 

`ifdef i_axi_AXI_R7_NEA_S16
  `define AXI_R7_NEA_S16 `i_axi_AXI_R7_NEA_S16
`endif 

`ifdef i_axi_AXI_R8_NSA_S1
  `define AXI_R8_NSA_S1 `i_axi_AXI_R8_NSA_S1
`endif 

`ifdef i_axi_AXI_R8_NEA_S1
  `define AXI_R8_NEA_S1 `i_axi_AXI_R8_NEA_S1
`endif 

`ifdef i_axi_AXI_R8_NSA_S2
  `define AXI_R8_NSA_S2 `i_axi_AXI_R8_NSA_S2
`endif 

`ifdef i_axi_AXI_R8_NEA_S2
  `define AXI_R8_NEA_S2 `i_axi_AXI_R8_NEA_S2
`endif 

`ifdef i_axi_AXI_R8_NSA_S3
  `define AXI_R8_NSA_S3 `i_axi_AXI_R8_NSA_S3
`endif 

`ifdef i_axi_AXI_R8_NEA_S3
  `define AXI_R8_NEA_S3 `i_axi_AXI_R8_NEA_S3
`endif 

`ifdef i_axi_AXI_R8_NSA_S4
  `define AXI_R8_NSA_S4 `i_axi_AXI_R8_NSA_S4
`endif 

`ifdef i_axi_AXI_R8_NEA_S4
  `define AXI_R8_NEA_S4 `i_axi_AXI_R8_NEA_S4
`endif 

`ifdef i_axi_AXI_R8_NSA_S5
  `define AXI_R8_NSA_S5 `i_axi_AXI_R8_NSA_S5
`endif 

`ifdef i_axi_AXI_R8_NEA_S5
  `define AXI_R8_NEA_S5 `i_axi_AXI_R8_NEA_S5
`endif 

`ifdef i_axi_AXI_R8_NSA_S6
  `define AXI_R8_NSA_S6 `i_axi_AXI_R8_NSA_S6
`endif 

`ifdef i_axi_AXI_R8_NEA_S6
  `define AXI_R8_NEA_S6 `i_axi_AXI_R8_NEA_S6
`endif 

`ifdef i_axi_AXI_R8_NSA_S7
  `define AXI_R8_NSA_S7 `i_axi_AXI_R8_NSA_S7
`endif 

`ifdef i_axi_AXI_R8_NEA_S7
  `define AXI_R8_NEA_S7 `i_axi_AXI_R8_NEA_S7
`endif 

`ifdef i_axi_AXI_R8_NSA_S8
  `define AXI_R8_NSA_S8 `i_axi_AXI_R8_NSA_S8
`endif 

`ifdef i_axi_AXI_R8_NEA_S8
  `define AXI_R8_NEA_S8 `i_axi_AXI_R8_NEA_S8
`endif 

`ifdef i_axi_AXI_R8_NSA_S9
  `define AXI_R8_NSA_S9 `i_axi_AXI_R8_NSA_S9
`endif 

`ifdef i_axi_AXI_R8_NEA_S9
  `define AXI_R8_NEA_S9 `i_axi_AXI_R8_NEA_S9
`endif 

`ifdef i_axi_AXI_R8_NSA_S10
  `define AXI_R8_NSA_S10 `i_axi_AXI_R8_NSA_S10
`endif 

`ifdef i_axi_AXI_R8_NEA_S10
  `define AXI_R8_NEA_S10 `i_axi_AXI_R8_NEA_S10
`endif 

`ifdef i_axi_AXI_R8_NSA_S11
  `define AXI_R8_NSA_S11 `i_axi_AXI_R8_NSA_S11
`endif 

`ifdef i_axi_AXI_R8_NEA_S11
  `define AXI_R8_NEA_S11 `i_axi_AXI_R8_NEA_S11
`endif 

`ifdef i_axi_AXI_R8_NSA_S12
  `define AXI_R8_NSA_S12 `i_axi_AXI_R8_NSA_S12
`endif 

`ifdef i_axi_AXI_R8_NEA_S12
  `define AXI_R8_NEA_S12 `i_axi_AXI_R8_NEA_S12
`endif 

`ifdef i_axi_AXI_R8_NSA_S13
  `define AXI_R8_NSA_S13 `i_axi_AXI_R8_NSA_S13
`endif 

`ifdef i_axi_AXI_R8_NEA_S13
  `define AXI_R8_NEA_S13 `i_axi_AXI_R8_NEA_S13
`endif 

`ifdef i_axi_AXI_R8_NSA_S14
  `define AXI_R8_NSA_S14 `i_axi_AXI_R8_NSA_S14
`endif 

`ifdef i_axi_AXI_R8_NEA_S14
  `define AXI_R8_NEA_S14 `i_axi_AXI_R8_NEA_S14
`endif 

`ifdef i_axi_AXI_R8_NSA_S15
  `define AXI_R8_NSA_S15 `i_axi_AXI_R8_NSA_S15
`endif 

`ifdef i_axi_AXI_R8_NEA_S15
  `define AXI_R8_NEA_S15 `i_axi_AXI_R8_NEA_S15
`endif 

`ifdef i_axi_AXI_R8_NSA_S16
  `define AXI_R8_NSA_S16 `i_axi_AXI_R8_NSA_S16
`endif 

`ifdef i_axi_AXI_R8_NEA_S16
  `define AXI_R8_NEA_S16 `i_axi_AXI_R8_NEA_S16
`endif 

`ifdef i_axi_AXI_NUM_RB_S1
  `define AXI_NUM_RB_S1 `i_axi_AXI_NUM_RB_S1
`endif 

`ifdef i_axi_AXI_NUM_RB_S2
  `define AXI_NUM_RB_S2 `i_axi_AXI_NUM_RB_S2
`endif 

`ifdef i_axi_AXI_NUM_RB_S3
  `define AXI_NUM_RB_S3 `i_axi_AXI_NUM_RB_S3
`endif 

`ifdef i_axi_AXI_NUM_RB_S4
  `define AXI_NUM_RB_S4 `i_axi_AXI_NUM_RB_S4
`endif 

`ifdef i_axi_AXI_NUM_RB_S5
  `define AXI_NUM_RB_S5 `i_axi_AXI_NUM_RB_S5
`endif 

`ifdef i_axi_AXI_NUM_RB_S6
  `define AXI_NUM_RB_S6 `i_axi_AXI_NUM_RB_S6
`endif 

`ifdef i_axi_AXI_NUM_RB_S7
  `define AXI_NUM_RB_S7 `i_axi_AXI_NUM_RB_S7
`endif 

`ifdef i_axi_AXI_NUM_RB_S8
  `define AXI_NUM_RB_S8 `i_axi_AXI_NUM_RB_S8
`endif 

`ifdef i_axi_AXI_NUM_RB_S9
  `define AXI_NUM_RB_S9 `i_axi_AXI_NUM_RB_S9
`endif 

`ifdef i_axi_AXI_NUM_RB_S10
  `define AXI_NUM_RB_S10 `i_axi_AXI_NUM_RB_S10
`endif 

`ifdef i_axi_AXI_NUM_RB_S11
  `define AXI_NUM_RB_S11 `i_axi_AXI_NUM_RB_S11
`endif 

`ifdef i_axi_AXI_NUM_RB_S12
  `define AXI_NUM_RB_S12 `i_axi_AXI_NUM_RB_S12
`endif 

`ifdef i_axi_AXI_NUM_RB_S13
  `define AXI_NUM_RB_S13 `i_axi_AXI_NUM_RB_S13
`endif 

`ifdef i_axi_AXI_NUM_RB_S14
  `define AXI_NUM_RB_S14 `i_axi_AXI_NUM_RB_S14
`endif 

`ifdef i_axi_AXI_NUM_RB_S15
  `define AXI_NUM_RB_S15 `i_axi_AXI_NUM_RB_S15
`endif 

`ifdef i_axi_AXI_NUM_RB_S16
  `define AXI_NUM_RB_S16 `i_axi_AXI_NUM_RB_S16
`endif 

`ifdef i_axi_AXI_R1_BSA_S1
  `define AXI_R1_BSA_S1 `i_axi_AXI_R1_BSA_S1
`endif 

`ifdef i_axi_AXI_R1_BEA_S1
  `define AXI_R1_BEA_S1 `i_axi_AXI_R1_BEA_S1
`endif 

`ifdef i_axi_AXI_R1_BSA_S2
  `define AXI_R1_BSA_S2 `i_axi_AXI_R1_BSA_S2
`endif 

`ifdef i_axi_AXI_R1_BEA_S2
  `define AXI_R1_BEA_S2 `i_axi_AXI_R1_BEA_S2
`endif 

`ifdef i_axi_AXI_R1_BSA_S3
  `define AXI_R1_BSA_S3 `i_axi_AXI_R1_BSA_S3
`endif 

`ifdef i_axi_AXI_R1_BEA_S3
  `define AXI_R1_BEA_S3 `i_axi_AXI_R1_BEA_S3
`endif 

`ifdef i_axi_AXI_R1_BSA_S4
  `define AXI_R1_BSA_S4 `i_axi_AXI_R1_BSA_S4
`endif 

`ifdef i_axi_AXI_R1_BEA_S4
  `define AXI_R1_BEA_S4 `i_axi_AXI_R1_BEA_S4
`endif 

`ifdef i_axi_AXI_R1_BSA_S5
  `define AXI_R1_BSA_S5 `i_axi_AXI_R1_BSA_S5
`endif 

`ifdef i_axi_AXI_R1_BEA_S5
  `define AXI_R1_BEA_S5 `i_axi_AXI_R1_BEA_S5
`endif 

`ifdef i_axi_AXI_R1_BSA_S6
  `define AXI_R1_BSA_S6 `i_axi_AXI_R1_BSA_S6
`endif 

`ifdef i_axi_AXI_R1_BEA_S6
  `define AXI_R1_BEA_S6 `i_axi_AXI_R1_BEA_S6
`endif 

`ifdef i_axi_AXI_R1_BSA_S7
  `define AXI_R1_BSA_S7 `i_axi_AXI_R1_BSA_S7
`endif 

`ifdef i_axi_AXI_R1_BEA_S7
  `define AXI_R1_BEA_S7 `i_axi_AXI_R1_BEA_S7
`endif 

`ifdef i_axi_AXI_R1_BSA_S8
  `define AXI_R1_BSA_S8 `i_axi_AXI_R1_BSA_S8
`endif 

`ifdef i_axi_AXI_R1_BEA_S8
  `define AXI_R1_BEA_S8 `i_axi_AXI_R1_BEA_S8
`endif 

`ifdef i_axi_AXI_R1_BSA_S9
  `define AXI_R1_BSA_S9 `i_axi_AXI_R1_BSA_S9
`endif 

`ifdef i_axi_AXI_R1_BEA_S9
  `define AXI_R1_BEA_S9 `i_axi_AXI_R1_BEA_S9
`endif 

`ifdef i_axi_AXI_R1_BSA_S10
  `define AXI_R1_BSA_S10 `i_axi_AXI_R1_BSA_S10
`endif 

`ifdef i_axi_AXI_R1_BEA_S10
  `define AXI_R1_BEA_S10 `i_axi_AXI_R1_BEA_S10
`endif 

`ifdef i_axi_AXI_R1_BSA_S11
  `define AXI_R1_BSA_S11 `i_axi_AXI_R1_BSA_S11
`endif 

`ifdef i_axi_AXI_R1_BEA_S11
  `define AXI_R1_BEA_S11 `i_axi_AXI_R1_BEA_S11
`endif 

`ifdef i_axi_AXI_R1_BSA_S12
  `define AXI_R1_BSA_S12 `i_axi_AXI_R1_BSA_S12
`endif 

`ifdef i_axi_AXI_R1_BEA_S12
  `define AXI_R1_BEA_S12 `i_axi_AXI_R1_BEA_S12
`endif 

`ifdef i_axi_AXI_R1_BSA_S13
  `define AXI_R1_BSA_S13 `i_axi_AXI_R1_BSA_S13
`endif 

`ifdef i_axi_AXI_R1_BEA_S13
  `define AXI_R1_BEA_S13 `i_axi_AXI_R1_BEA_S13
`endif 

`ifdef i_axi_AXI_R1_BSA_S14
  `define AXI_R1_BSA_S14 `i_axi_AXI_R1_BSA_S14
`endif 

`ifdef i_axi_AXI_R1_BEA_S14
  `define AXI_R1_BEA_S14 `i_axi_AXI_R1_BEA_S14
`endif 

`ifdef i_axi_AXI_R1_BSA_S15
  `define AXI_R1_BSA_S15 `i_axi_AXI_R1_BSA_S15
`endif 

`ifdef i_axi_AXI_R1_BEA_S15
  `define AXI_R1_BEA_S15 `i_axi_AXI_R1_BEA_S15
`endif 

`ifdef i_axi_AXI_R1_BSA_S16
  `define AXI_R1_BSA_S16 `i_axi_AXI_R1_BSA_S16
`endif 

`ifdef i_axi_AXI_R1_BEA_S16
  `define AXI_R1_BEA_S16 `i_axi_AXI_R1_BEA_S16
`endif 

`ifdef i_axi_AXI_R2_BSA_S1
  `define AXI_R2_BSA_S1 `i_axi_AXI_R2_BSA_S1
`endif 

`ifdef i_axi_AXI_R2_BEA_S1
  `define AXI_R2_BEA_S1 `i_axi_AXI_R2_BEA_S1
`endif 

`ifdef i_axi_AXI_R2_BSA_S2
  `define AXI_R2_BSA_S2 `i_axi_AXI_R2_BSA_S2
`endif 

`ifdef i_axi_AXI_R2_BEA_S2
  `define AXI_R2_BEA_S2 `i_axi_AXI_R2_BEA_S2
`endif 

`ifdef i_axi_AXI_R2_BSA_S3
  `define AXI_R2_BSA_S3 `i_axi_AXI_R2_BSA_S3
`endif 

`ifdef i_axi_AXI_R2_BEA_S3
  `define AXI_R2_BEA_S3 `i_axi_AXI_R2_BEA_S3
`endif 

`ifdef i_axi_AXI_R2_BSA_S4
  `define AXI_R2_BSA_S4 `i_axi_AXI_R2_BSA_S4
`endif 

`ifdef i_axi_AXI_R2_BEA_S4
  `define AXI_R2_BEA_S4 `i_axi_AXI_R2_BEA_S4
`endif 

`ifdef i_axi_AXI_R2_BSA_S5
  `define AXI_R2_BSA_S5 `i_axi_AXI_R2_BSA_S5
`endif 

`ifdef i_axi_AXI_R2_BEA_S5
  `define AXI_R2_BEA_S5 `i_axi_AXI_R2_BEA_S5
`endif 

`ifdef i_axi_AXI_R2_BSA_S6
  `define AXI_R2_BSA_S6 `i_axi_AXI_R2_BSA_S6
`endif 

`ifdef i_axi_AXI_R2_BEA_S6
  `define AXI_R2_BEA_S6 `i_axi_AXI_R2_BEA_S6
`endif 

`ifdef i_axi_AXI_R2_BSA_S7
  `define AXI_R2_BSA_S7 `i_axi_AXI_R2_BSA_S7
`endif 

`ifdef i_axi_AXI_R2_BEA_S7
  `define AXI_R2_BEA_S7 `i_axi_AXI_R2_BEA_S7
`endif 

`ifdef i_axi_AXI_R2_BSA_S8
  `define AXI_R2_BSA_S8 `i_axi_AXI_R2_BSA_S8
`endif 

`ifdef i_axi_AXI_R2_BEA_S8
  `define AXI_R2_BEA_S8 `i_axi_AXI_R2_BEA_S8
`endif 

`ifdef i_axi_AXI_R2_BSA_S9
  `define AXI_R2_BSA_S9 `i_axi_AXI_R2_BSA_S9
`endif 

`ifdef i_axi_AXI_R2_BEA_S9
  `define AXI_R2_BEA_S9 `i_axi_AXI_R2_BEA_S9
`endif 

`ifdef i_axi_AXI_R2_BSA_S10
  `define AXI_R2_BSA_S10 `i_axi_AXI_R2_BSA_S10
`endif 

`ifdef i_axi_AXI_R2_BEA_S10
  `define AXI_R2_BEA_S10 `i_axi_AXI_R2_BEA_S10
`endif 

`ifdef i_axi_AXI_R2_BSA_S11
  `define AXI_R2_BSA_S11 `i_axi_AXI_R2_BSA_S11
`endif 

`ifdef i_axi_AXI_R2_BEA_S11
  `define AXI_R2_BEA_S11 `i_axi_AXI_R2_BEA_S11
`endif 

`ifdef i_axi_AXI_R2_BSA_S12
  `define AXI_R2_BSA_S12 `i_axi_AXI_R2_BSA_S12
`endif 

`ifdef i_axi_AXI_R2_BEA_S12
  `define AXI_R2_BEA_S12 `i_axi_AXI_R2_BEA_S12
`endif 

`ifdef i_axi_AXI_R2_BSA_S13
  `define AXI_R2_BSA_S13 `i_axi_AXI_R2_BSA_S13
`endif 

`ifdef i_axi_AXI_R2_BEA_S13
  `define AXI_R2_BEA_S13 `i_axi_AXI_R2_BEA_S13
`endif 

`ifdef i_axi_AXI_R2_BSA_S14
  `define AXI_R2_BSA_S14 `i_axi_AXI_R2_BSA_S14
`endif 

`ifdef i_axi_AXI_R2_BEA_S14
  `define AXI_R2_BEA_S14 `i_axi_AXI_R2_BEA_S14
`endif 

`ifdef i_axi_AXI_R2_BSA_S15
  `define AXI_R2_BSA_S15 `i_axi_AXI_R2_BSA_S15
`endif 

`ifdef i_axi_AXI_R2_BEA_S15
  `define AXI_R2_BEA_S15 `i_axi_AXI_R2_BEA_S15
`endif 

`ifdef i_axi_AXI_R2_BSA_S16
  `define AXI_R2_BSA_S16 `i_axi_AXI_R2_BSA_S16
`endif 

`ifdef i_axi_AXI_R2_BEA_S16
  `define AXI_R2_BEA_S16 `i_axi_AXI_R2_BEA_S16
`endif 

`ifdef i_axi_AXI_R3_BSA_S1
  `define AXI_R3_BSA_S1 `i_axi_AXI_R3_BSA_S1
`endif 

`ifdef i_axi_AXI_R3_BEA_S1
  `define AXI_R3_BEA_S1 `i_axi_AXI_R3_BEA_S1
`endif 

`ifdef i_axi_AXI_R3_BSA_S2
  `define AXI_R3_BSA_S2 `i_axi_AXI_R3_BSA_S2
`endif 

`ifdef i_axi_AXI_R3_BEA_S2
  `define AXI_R3_BEA_S2 `i_axi_AXI_R3_BEA_S2
`endif 

`ifdef i_axi_AXI_R3_BSA_S3
  `define AXI_R3_BSA_S3 `i_axi_AXI_R3_BSA_S3
`endif 

`ifdef i_axi_AXI_R3_BEA_S3
  `define AXI_R3_BEA_S3 `i_axi_AXI_R3_BEA_S3
`endif 

`ifdef i_axi_AXI_R3_BSA_S4
  `define AXI_R3_BSA_S4 `i_axi_AXI_R3_BSA_S4
`endif 

`ifdef i_axi_AXI_R3_BEA_S4
  `define AXI_R3_BEA_S4 `i_axi_AXI_R3_BEA_S4
`endif 

`ifdef i_axi_AXI_R3_BSA_S5
  `define AXI_R3_BSA_S5 `i_axi_AXI_R3_BSA_S5
`endif 

`ifdef i_axi_AXI_R3_BEA_S5
  `define AXI_R3_BEA_S5 `i_axi_AXI_R3_BEA_S5
`endif 

`ifdef i_axi_AXI_R3_BSA_S6
  `define AXI_R3_BSA_S6 `i_axi_AXI_R3_BSA_S6
`endif 

`ifdef i_axi_AXI_R3_BEA_S6
  `define AXI_R3_BEA_S6 `i_axi_AXI_R3_BEA_S6
`endif 

`ifdef i_axi_AXI_R3_BSA_S7
  `define AXI_R3_BSA_S7 `i_axi_AXI_R3_BSA_S7
`endif 

`ifdef i_axi_AXI_R3_BEA_S7
  `define AXI_R3_BEA_S7 `i_axi_AXI_R3_BEA_S7
`endif 

`ifdef i_axi_AXI_R3_BSA_S8
  `define AXI_R3_BSA_S8 `i_axi_AXI_R3_BSA_S8
`endif 

`ifdef i_axi_AXI_R3_BEA_S8
  `define AXI_R3_BEA_S8 `i_axi_AXI_R3_BEA_S8
`endif 

`ifdef i_axi_AXI_R3_BSA_S9
  `define AXI_R3_BSA_S9 `i_axi_AXI_R3_BSA_S9
`endif 

`ifdef i_axi_AXI_R3_BEA_S9
  `define AXI_R3_BEA_S9 `i_axi_AXI_R3_BEA_S9
`endif 

`ifdef i_axi_AXI_R3_BSA_S10
  `define AXI_R3_BSA_S10 `i_axi_AXI_R3_BSA_S10
`endif 

`ifdef i_axi_AXI_R3_BEA_S10
  `define AXI_R3_BEA_S10 `i_axi_AXI_R3_BEA_S10
`endif 

`ifdef i_axi_AXI_R3_BSA_S11
  `define AXI_R3_BSA_S11 `i_axi_AXI_R3_BSA_S11
`endif 

`ifdef i_axi_AXI_R3_BEA_S11
  `define AXI_R3_BEA_S11 `i_axi_AXI_R3_BEA_S11
`endif 

`ifdef i_axi_AXI_R3_BSA_S12
  `define AXI_R3_BSA_S12 `i_axi_AXI_R3_BSA_S12
`endif 

`ifdef i_axi_AXI_R3_BEA_S12
  `define AXI_R3_BEA_S12 `i_axi_AXI_R3_BEA_S12
`endif 

`ifdef i_axi_AXI_R3_BSA_S13
  `define AXI_R3_BSA_S13 `i_axi_AXI_R3_BSA_S13
`endif 

`ifdef i_axi_AXI_R3_BEA_S13
  `define AXI_R3_BEA_S13 `i_axi_AXI_R3_BEA_S13
`endif 

`ifdef i_axi_AXI_R3_BSA_S14
  `define AXI_R3_BSA_S14 `i_axi_AXI_R3_BSA_S14
`endif 

`ifdef i_axi_AXI_R3_BEA_S14
  `define AXI_R3_BEA_S14 `i_axi_AXI_R3_BEA_S14
`endif 

`ifdef i_axi_AXI_R3_BSA_S15
  `define AXI_R3_BSA_S15 `i_axi_AXI_R3_BSA_S15
`endif 

`ifdef i_axi_AXI_R3_BEA_S15
  `define AXI_R3_BEA_S15 `i_axi_AXI_R3_BEA_S15
`endif 

`ifdef i_axi_AXI_R3_BSA_S16
  `define AXI_R3_BSA_S16 `i_axi_AXI_R3_BSA_S16
`endif 

`ifdef i_axi_AXI_R3_BEA_S16
  `define AXI_R3_BEA_S16 `i_axi_AXI_R3_BEA_S16
`endif 

`ifdef i_axi_AXI_R4_BSA_S1
  `define AXI_R4_BSA_S1 `i_axi_AXI_R4_BSA_S1
`endif 

`ifdef i_axi_AXI_R4_BEA_S1
  `define AXI_R4_BEA_S1 `i_axi_AXI_R4_BEA_S1
`endif 

`ifdef i_axi_AXI_R4_BSA_S2
  `define AXI_R4_BSA_S2 `i_axi_AXI_R4_BSA_S2
`endif 

`ifdef i_axi_AXI_R4_BEA_S2
  `define AXI_R4_BEA_S2 `i_axi_AXI_R4_BEA_S2
`endif 

`ifdef i_axi_AXI_R4_BSA_S3
  `define AXI_R4_BSA_S3 `i_axi_AXI_R4_BSA_S3
`endif 

`ifdef i_axi_AXI_R4_BEA_S3
  `define AXI_R4_BEA_S3 `i_axi_AXI_R4_BEA_S3
`endif 

`ifdef i_axi_AXI_R4_BSA_S4
  `define AXI_R4_BSA_S4 `i_axi_AXI_R4_BSA_S4
`endif 

`ifdef i_axi_AXI_R4_BEA_S4
  `define AXI_R4_BEA_S4 `i_axi_AXI_R4_BEA_S4
`endif 

`ifdef i_axi_AXI_R4_BSA_S5
  `define AXI_R4_BSA_S5 `i_axi_AXI_R4_BSA_S5
`endif 

`ifdef i_axi_AXI_R4_BEA_S5
  `define AXI_R4_BEA_S5 `i_axi_AXI_R4_BEA_S5
`endif 

`ifdef i_axi_AXI_R4_BSA_S6
  `define AXI_R4_BSA_S6 `i_axi_AXI_R4_BSA_S6
`endif 

`ifdef i_axi_AXI_R4_BEA_S6
  `define AXI_R4_BEA_S6 `i_axi_AXI_R4_BEA_S6
`endif 

`ifdef i_axi_AXI_R4_BSA_S7
  `define AXI_R4_BSA_S7 `i_axi_AXI_R4_BSA_S7
`endif 

`ifdef i_axi_AXI_R4_BEA_S7
  `define AXI_R4_BEA_S7 `i_axi_AXI_R4_BEA_S7
`endif 

`ifdef i_axi_AXI_R4_BSA_S8
  `define AXI_R4_BSA_S8 `i_axi_AXI_R4_BSA_S8
`endif 

`ifdef i_axi_AXI_R4_BEA_S8
  `define AXI_R4_BEA_S8 `i_axi_AXI_R4_BEA_S8
`endif 

`ifdef i_axi_AXI_R4_BSA_S9
  `define AXI_R4_BSA_S9 `i_axi_AXI_R4_BSA_S9
`endif 

`ifdef i_axi_AXI_R4_BEA_S9
  `define AXI_R4_BEA_S9 `i_axi_AXI_R4_BEA_S9
`endif 

`ifdef i_axi_AXI_R4_BSA_S10
  `define AXI_R4_BSA_S10 `i_axi_AXI_R4_BSA_S10
`endif 

`ifdef i_axi_AXI_R4_BEA_S10
  `define AXI_R4_BEA_S10 `i_axi_AXI_R4_BEA_S10
`endif 

`ifdef i_axi_AXI_R4_BSA_S11
  `define AXI_R4_BSA_S11 `i_axi_AXI_R4_BSA_S11
`endif 

`ifdef i_axi_AXI_R4_BEA_S11
  `define AXI_R4_BEA_S11 `i_axi_AXI_R4_BEA_S11
`endif 

`ifdef i_axi_AXI_R4_BSA_S12
  `define AXI_R4_BSA_S12 `i_axi_AXI_R4_BSA_S12
`endif 

`ifdef i_axi_AXI_R4_BEA_S12
  `define AXI_R4_BEA_S12 `i_axi_AXI_R4_BEA_S12
`endif 

`ifdef i_axi_AXI_R4_BSA_S13
  `define AXI_R4_BSA_S13 `i_axi_AXI_R4_BSA_S13
`endif 

`ifdef i_axi_AXI_R4_BEA_S13
  `define AXI_R4_BEA_S13 `i_axi_AXI_R4_BEA_S13
`endif 

`ifdef i_axi_AXI_R4_BSA_S14
  `define AXI_R4_BSA_S14 `i_axi_AXI_R4_BSA_S14
`endif 

`ifdef i_axi_AXI_R4_BEA_S14
  `define AXI_R4_BEA_S14 `i_axi_AXI_R4_BEA_S14
`endif 

`ifdef i_axi_AXI_R4_BSA_S15
  `define AXI_R4_BSA_S15 `i_axi_AXI_R4_BSA_S15
`endif 

`ifdef i_axi_AXI_R4_BEA_S15
  `define AXI_R4_BEA_S15 `i_axi_AXI_R4_BEA_S15
`endif 

`ifdef i_axi_AXI_R4_BSA_S16
  `define AXI_R4_BSA_S16 `i_axi_AXI_R4_BSA_S16
`endif 

`ifdef i_axi_AXI_R4_BEA_S16
  `define AXI_R4_BEA_S16 `i_axi_AXI_R4_BEA_S16
`endif 

`ifdef i_axi_AXI_R5_BSA_S1
  `define AXI_R5_BSA_S1 `i_axi_AXI_R5_BSA_S1
`endif 

`ifdef i_axi_AXI_R5_BEA_S1
  `define AXI_R5_BEA_S1 `i_axi_AXI_R5_BEA_S1
`endif 

`ifdef i_axi_AXI_R5_BSA_S2
  `define AXI_R5_BSA_S2 `i_axi_AXI_R5_BSA_S2
`endif 

`ifdef i_axi_AXI_R5_BEA_S2
  `define AXI_R5_BEA_S2 `i_axi_AXI_R5_BEA_S2
`endif 

`ifdef i_axi_AXI_R5_BSA_S3
  `define AXI_R5_BSA_S3 `i_axi_AXI_R5_BSA_S3
`endif 

`ifdef i_axi_AXI_R5_BEA_S3
  `define AXI_R5_BEA_S3 `i_axi_AXI_R5_BEA_S3
`endif 

`ifdef i_axi_AXI_R5_BSA_S4
  `define AXI_R5_BSA_S4 `i_axi_AXI_R5_BSA_S4
`endif 

`ifdef i_axi_AXI_R5_BEA_S4
  `define AXI_R5_BEA_S4 `i_axi_AXI_R5_BEA_S4
`endif 

`ifdef i_axi_AXI_R5_BSA_S5
  `define AXI_R5_BSA_S5 `i_axi_AXI_R5_BSA_S5
`endif 

`ifdef i_axi_AXI_R5_BEA_S5
  `define AXI_R5_BEA_S5 `i_axi_AXI_R5_BEA_S5
`endif 

`ifdef i_axi_AXI_R5_BSA_S6
  `define AXI_R5_BSA_S6 `i_axi_AXI_R5_BSA_S6
`endif 

`ifdef i_axi_AXI_R5_BEA_S6
  `define AXI_R5_BEA_S6 `i_axi_AXI_R5_BEA_S6
`endif 

`ifdef i_axi_AXI_R5_BSA_S7
  `define AXI_R5_BSA_S7 `i_axi_AXI_R5_BSA_S7
`endif 

`ifdef i_axi_AXI_R5_BEA_S7
  `define AXI_R5_BEA_S7 `i_axi_AXI_R5_BEA_S7
`endif 

`ifdef i_axi_AXI_R5_BSA_S8
  `define AXI_R5_BSA_S8 `i_axi_AXI_R5_BSA_S8
`endif 

`ifdef i_axi_AXI_R5_BEA_S8
  `define AXI_R5_BEA_S8 `i_axi_AXI_R5_BEA_S8
`endif 

`ifdef i_axi_AXI_R5_BSA_S9
  `define AXI_R5_BSA_S9 `i_axi_AXI_R5_BSA_S9
`endif 

`ifdef i_axi_AXI_R5_BEA_S9
  `define AXI_R5_BEA_S9 `i_axi_AXI_R5_BEA_S9
`endif 

`ifdef i_axi_AXI_R5_BSA_S10
  `define AXI_R5_BSA_S10 `i_axi_AXI_R5_BSA_S10
`endif 

`ifdef i_axi_AXI_R5_BEA_S10
  `define AXI_R5_BEA_S10 `i_axi_AXI_R5_BEA_S10
`endif 

`ifdef i_axi_AXI_R5_BSA_S11
  `define AXI_R5_BSA_S11 `i_axi_AXI_R5_BSA_S11
`endif 

`ifdef i_axi_AXI_R5_BEA_S11
  `define AXI_R5_BEA_S11 `i_axi_AXI_R5_BEA_S11
`endif 

`ifdef i_axi_AXI_R5_BSA_S12
  `define AXI_R5_BSA_S12 `i_axi_AXI_R5_BSA_S12
`endif 

`ifdef i_axi_AXI_R5_BEA_S12
  `define AXI_R5_BEA_S12 `i_axi_AXI_R5_BEA_S12
`endif 

`ifdef i_axi_AXI_R5_BSA_S13
  `define AXI_R5_BSA_S13 `i_axi_AXI_R5_BSA_S13
`endif 

`ifdef i_axi_AXI_R5_BEA_S13
  `define AXI_R5_BEA_S13 `i_axi_AXI_R5_BEA_S13
`endif 

`ifdef i_axi_AXI_R5_BSA_S14
  `define AXI_R5_BSA_S14 `i_axi_AXI_R5_BSA_S14
`endif 

`ifdef i_axi_AXI_R5_BEA_S14
  `define AXI_R5_BEA_S14 `i_axi_AXI_R5_BEA_S14
`endif 

`ifdef i_axi_AXI_R5_BSA_S15
  `define AXI_R5_BSA_S15 `i_axi_AXI_R5_BSA_S15
`endif 

`ifdef i_axi_AXI_R5_BEA_S15
  `define AXI_R5_BEA_S15 `i_axi_AXI_R5_BEA_S15
`endif 

`ifdef i_axi_AXI_R5_BSA_S16
  `define AXI_R5_BSA_S16 `i_axi_AXI_R5_BSA_S16
`endif 

`ifdef i_axi_AXI_R5_BEA_S16
  `define AXI_R5_BEA_S16 `i_axi_AXI_R5_BEA_S16
`endif 

`ifdef i_axi_AXI_R6_BSA_S1
  `define AXI_R6_BSA_S1 `i_axi_AXI_R6_BSA_S1
`endif 

`ifdef i_axi_AXI_R6_BEA_S1
  `define AXI_R6_BEA_S1 `i_axi_AXI_R6_BEA_S1
`endif 

`ifdef i_axi_AXI_R6_BSA_S2
  `define AXI_R6_BSA_S2 `i_axi_AXI_R6_BSA_S2
`endif 

`ifdef i_axi_AXI_R6_BEA_S2
  `define AXI_R6_BEA_S2 `i_axi_AXI_R6_BEA_S2
`endif 

`ifdef i_axi_AXI_R6_BSA_S3
  `define AXI_R6_BSA_S3 `i_axi_AXI_R6_BSA_S3
`endif 

`ifdef i_axi_AXI_R6_BEA_S3
  `define AXI_R6_BEA_S3 `i_axi_AXI_R6_BEA_S3
`endif 

`ifdef i_axi_AXI_R6_BSA_S4
  `define AXI_R6_BSA_S4 `i_axi_AXI_R6_BSA_S4
`endif 

`ifdef i_axi_AXI_R6_BEA_S4
  `define AXI_R6_BEA_S4 `i_axi_AXI_R6_BEA_S4
`endif 

`ifdef i_axi_AXI_R6_BSA_S5
  `define AXI_R6_BSA_S5 `i_axi_AXI_R6_BSA_S5
`endif 

`ifdef i_axi_AXI_R6_BEA_S5
  `define AXI_R6_BEA_S5 `i_axi_AXI_R6_BEA_S5
`endif 

`ifdef i_axi_AXI_R6_BSA_S6
  `define AXI_R6_BSA_S6 `i_axi_AXI_R6_BSA_S6
`endif 

`ifdef i_axi_AXI_R6_BEA_S6
  `define AXI_R6_BEA_S6 `i_axi_AXI_R6_BEA_S6
`endif 

`ifdef i_axi_AXI_R6_BSA_S7
  `define AXI_R6_BSA_S7 `i_axi_AXI_R6_BSA_S7
`endif 

`ifdef i_axi_AXI_R6_BEA_S7
  `define AXI_R6_BEA_S7 `i_axi_AXI_R6_BEA_S7
`endif 

`ifdef i_axi_AXI_R6_BSA_S8
  `define AXI_R6_BSA_S8 `i_axi_AXI_R6_BSA_S8
`endif 

`ifdef i_axi_AXI_R6_BEA_S8
  `define AXI_R6_BEA_S8 `i_axi_AXI_R6_BEA_S8
`endif 

`ifdef i_axi_AXI_R6_BSA_S9
  `define AXI_R6_BSA_S9 `i_axi_AXI_R6_BSA_S9
`endif 

`ifdef i_axi_AXI_R6_BEA_S9
  `define AXI_R6_BEA_S9 `i_axi_AXI_R6_BEA_S9
`endif 

`ifdef i_axi_AXI_R6_BSA_S10
  `define AXI_R6_BSA_S10 `i_axi_AXI_R6_BSA_S10
`endif 

`ifdef i_axi_AXI_R6_BEA_S10
  `define AXI_R6_BEA_S10 `i_axi_AXI_R6_BEA_S10
`endif 

`ifdef i_axi_AXI_R6_BSA_S11
  `define AXI_R6_BSA_S11 `i_axi_AXI_R6_BSA_S11
`endif 

`ifdef i_axi_AXI_R6_BEA_S11
  `define AXI_R6_BEA_S11 `i_axi_AXI_R6_BEA_S11
`endif 

`ifdef i_axi_AXI_R6_BSA_S12
  `define AXI_R6_BSA_S12 `i_axi_AXI_R6_BSA_S12
`endif 

`ifdef i_axi_AXI_R6_BEA_S12
  `define AXI_R6_BEA_S12 `i_axi_AXI_R6_BEA_S12
`endif 

`ifdef i_axi_AXI_R6_BSA_S13
  `define AXI_R6_BSA_S13 `i_axi_AXI_R6_BSA_S13
`endif 

`ifdef i_axi_AXI_R6_BEA_S13
  `define AXI_R6_BEA_S13 `i_axi_AXI_R6_BEA_S13
`endif 

`ifdef i_axi_AXI_R6_BSA_S14
  `define AXI_R6_BSA_S14 `i_axi_AXI_R6_BSA_S14
`endif 

`ifdef i_axi_AXI_R6_BEA_S14
  `define AXI_R6_BEA_S14 `i_axi_AXI_R6_BEA_S14
`endif 

`ifdef i_axi_AXI_R6_BSA_S15
  `define AXI_R6_BSA_S15 `i_axi_AXI_R6_BSA_S15
`endif 

`ifdef i_axi_AXI_R6_BEA_S15
  `define AXI_R6_BEA_S15 `i_axi_AXI_R6_BEA_S15
`endif 

`ifdef i_axi_AXI_R6_BSA_S16
  `define AXI_R6_BSA_S16 `i_axi_AXI_R6_BSA_S16
`endif 

`ifdef i_axi_AXI_R6_BEA_S16
  `define AXI_R6_BEA_S16 `i_axi_AXI_R6_BEA_S16
`endif 

`ifdef i_axi_AXI_R7_BSA_S1
  `define AXI_R7_BSA_S1 `i_axi_AXI_R7_BSA_S1
`endif 

`ifdef i_axi_AXI_R7_BEA_S1
  `define AXI_R7_BEA_S1 `i_axi_AXI_R7_BEA_S1
`endif 

`ifdef i_axi_AXI_R7_BSA_S2
  `define AXI_R7_BSA_S2 `i_axi_AXI_R7_BSA_S2
`endif 

`ifdef i_axi_AXI_R7_BEA_S2
  `define AXI_R7_BEA_S2 `i_axi_AXI_R7_BEA_S2
`endif 

`ifdef i_axi_AXI_R7_BSA_S3
  `define AXI_R7_BSA_S3 `i_axi_AXI_R7_BSA_S3
`endif 

`ifdef i_axi_AXI_R7_BEA_S3
  `define AXI_R7_BEA_S3 `i_axi_AXI_R7_BEA_S3
`endif 

`ifdef i_axi_AXI_R7_BSA_S4
  `define AXI_R7_BSA_S4 `i_axi_AXI_R7_BSA_S4
`endif 

`ifdef i_axi_AXI_R7_BEA_S4
  `define AXI_R7_BEA_S4 `i_axi_AXI_R7_BEA_S4
`endif 

`ifdef i_axi_AXI_R7_BSA_S5
  `define AXI_R7_BSA_S5 `i_axi_AXI_R7_BSA_S5
`endif 

`ifdef i_axi_AXI_R7_BEA_S5
  `define AXI_R7_BEA_S5 `i_axi_AXI_R7_BEA_S5
`endif 

`ifdef i_axi_AXI_R7_BSA_S6
  `define AXI_R7_BSA_S6 `i_axi_AXI_R7_BSA_S6
`endif 

`ifdef i_axi_AXI_R7_BEA_S6
  `define AXI_R7_BEA_S6 `i_axi_AXI_R7_BEA_S6
`endif 

`ifdef i_axi_AXI_R7_BSA_S7
  `define AXI_R7_BSA_S7 `i_axi_AXI_R7_BSA_S7
`endif 

`ifdef i_axi_AXI_R7_BEA_S7
  `define AXI_R7_BEA_S7 `i_axi_AXI_R7_BEA_S7
`endif 

`ifdef i_axi_AXI_R7_BSA_S8
  `define AXI_R7_BSA_S8 `i_axi_AXI_R7_BSA_S8
`endif 

`ifdef i_axi_AXI_R7_BEA_S8
  `define AXI_R7_BEA_S8 `i_axi_AXI_R7_BEA_S8
`endif 

`ifdef i_axi_AXI_R7_BSA_S9
  `define AXI_R7_BSA_S9 `i_axi_AXI_R7_BSA_S9
`endif 

`ifdef i_axi_AXI_R7_BEA_S9
  `define AXI_R7_BEA_S9 `i_axi_AXI_R7_BEA_S9
`endif 

`ifdef i_axi_AXI_R7_BSA_S10
  `define AXI_R7_BSA_S10 `i_axi_AXI_R7_BSA_S10
`endif 

`ifdef i_axi_AXI_R7_BEA_S10
  `define AXI_R7_BEA_S10 `i_axi_AXI_R7_BEA_S10
`endif 

`ifdef i_axi_AXI_R7_BSA_S11
  `define AXI_R7_BSA_S11 `i_axi_AXI_R7_BSA_S11
`endif 

`ifdef i_axi_AXI_R7_BEA_S11
  `define AXI_R7_BEA_S11 `i_axi_AXI_R7_BEA_S11
`endif 

`ifdef i_axi_AXI_R7_BSA_S12
  `define AXI_R7_BSA_S12 `i_axi_AXI_R7_BSA_S12
`endif 

`ifdef i_axi_AXI_R7_BEA_S12
  `define AXI_R7_BEA_S12 `i_axi_AXI_R7_BEA_S12
`endif 

`ifdef i_axi_AXI_R7_BSA_S13
  `define AXI_R7_BSA_S13 `i_axi_AXI_R7_BSA_S13
`endif 

`ifdef i_axi_AXI_R7_BEA_S13
  `define AXI_R7_BEA_S13 `i_axi_AXI_R7_BEA_S13
`endif 

`ifdef i_axi_AXI_R7_BSA_S14
  `define AXI_R7_BSA_S14 `i_axi_AXI_R7_BSA_S14
`endif 

`ifdef i_axi_AXI_R7_BEA_S14
  `define AXI_R7_BEA_S14 `i_axi_AXI_R7_BEA_S14
`endif 

`ifdef i_axi_AXI_R7_BSA_S15
  `define AXI_R7_BSA_S15 `i_axi_AXI_R7_BSA_S15
`endif 

`ifdef i_axi_AXI_R7_BEA_S15
  `define AXI_R7_BEA_S15 `i_axi_AXI_R7_BEA_S15
`endif 

`ifdef i_axi_AXI_R7_BSA_S16
  `define AXI_R7_BSA_S16 `i_axi_AXI_R7_BSA_S16
`endif 

`ifdef i_axi_AXI_R7_BEA_S16
  `define AXI_R7_BEA_S16 `i_axi_AXI_R7_BEA_S16
`endif 

`ifdef i_axi_AXI_R8_BSA_S1
  `define AXI_R8_BSA_S1 `i_axi_AXI_R8_BSA_S1
`endif 

`ifdef i_axi_AXI_R8_BEA_S1
  `define AXI_R8_BEA_S1 `i_axi_AXI_R8_BEA_S1
`endif 

`ifdef i_axi_AXI_R8_BSA_S2
  `define AXI_R8_BSA_S2 `i_axi_AXI_R8_BSA_S2
`endif 

`ifdef i_axi_AXI_R8_BEA_S2
  `define AXI_R8_BEA_S2 `i_axi_AXI_R8_BEA_S2
`endif 

`ifdef i_axi_AXI_R8_BSA_S3
  `define AXI_R8_BSA_S3 `i_axi_AXI_R8_BSA_S3
`endif 

`ifdef i_axi_AXI_R8_BEA_S3
  `define AXI_R8_BEA_S3 `i_axi_AXI_R8_BEA_S3
`endif 

`ifdef i_axi_AXI_R8_BSA_S4
  `define AXI_R8_BSA_S4 `i_axi_AXI_R8_BSA_S4
`endif 

`ifdef i_axi_AXI_R8_BEA_S4
  `define AXI_R8_BEA_S4 `i_axi_AXI_R8_BEA_S4
`endif 

`ifdef i_axi_AXI_R8_BSA_S5
  `define AXI_R8_BSA_S5 `i_axi_AXI_R8_BSA_S5
`endif 

`ifdef i_axi_AXI_R8_BEA_S5
  `define AXI_R8_BEA_S5 `i_axi_AXI_R8_BEA_S5
`endif 

`ifdef i_axi_AXI_R8_BSA_S6
  `define AXI_R8_BSA_S6 `i_axi_AXI_R8_BSA_S6
`endif 

`ifdef i_axi_AXI_R8_BEA_S6
  `define AXI_R8_BEA_S6 `i_axi_AXI_R8_BEA_S6
`endif 

`ifdef i_axi_AXI_R8_BSA_S7
  `define AXI_R8_BSA_S7 `i_axi_AXI_R8_BSA_S7
`endif 

`ifdef i_axi_AXI_R8_BEA_S7
  `define AXI_R8_BEA_S7 `i_axi_AXI_R8_BEA_S7
`endif 

`ifdef i_axi_AXI_R8_BSA_S8
  `define AXI_R8_BSA_S8 `i_axi_AXI_R8_BSA_S8
`endif 

`ifdef i_axi_AXI_R8_BEA_S8
  `define AXI_R8_BEA_S8 `i_axi_AXI_R8_BEA_S8
`endif 

`ifdef i_axi_AXI_R8_BSA_S9
  `define AXI_R8_BSA_S9 `i_axi_AXI_R8_BSA_S9
`endif 

`ifdef i_axi_AXI_R8_BEA_S9
  `define AXI_R8_BEA_S9 `i_axi_AXI_R8_BEA_S9
`endif 

`ifdef i_axi_AXI_R8_BSA_S10
  `define AXI_R8_BSA_S10 `i_axi_AXI_R8_BSA_S10
`endif 

`ifdef i_axi_AXI_R8_BEA_S10
  `define AXI_R8_BEA_S10 `i_axi_AXI_R8_BEA_S10
`endif 

`ifdef i_axi_AXI_R8_BSA_S11
  `define AXI_R8_BSA_S11 `i_axi_AXI_R8_BSA_S11
`endif 

`ifdef i_axi_AXI_R8_BEA_S11
  `define AXI_R8_BEA_S11 `i_axi_AXI_R8_BEA_S11
`endif 

`ifdef i_axi_AXI_R8_BSA_S12
  `define AXI_R8_BSA_S12 `i_axi_AXI_R8_BSA_S12
`endif 

`ifdef i_axi_AXI_R8_BEA_S12
  `define AXI_R8_BEA_S12 `i_axi_AXI_R8_BEA_S12
`endif 

`ifdef i_axi_AXI_R8_BSA_S13
  `define AXI_R8_BSA_S13 `i_axi_AXI_R8_BSA_S13
`endif 

`ifdef i_axi_AXI_R8_BEA_S13
  `define AXI_R8_BEA_S13 `i_axi_AXI_R8_BEA_S13
`endif 

`ifdef i_axi_AXI_R8_BSA_S14
  `define AXI_R8_BSA_S14 `i_axi_AXI_R8_BSA_S14
`endif 

`ifdef i_axi_AXI_R8_BEA_S14
  `define AXI_R8_BEA_S14 `i_axi_AXI_R8_BEA_S14
`endif 

`ifdef i_axi_AXI_R8_BSA_S15
  `define AXI_R8_BSA_S15 `i_axi_AXI_R8_BSA_S15
`endif 

`ifdef i_axi_AXI_R8_BEA_S15
  `define AXI_R8_BEA_S15 `i_axi_AXI_R8_BEA_S15
`endif 

`ifdef i_axi_AXI_R8_BSA_S16
  `define AXI_R8_BSA_S16 `i_axi_AXI_R8_BSA_S16
`endif 

`ifdef i_axi_AXI_R8_BEA_S16
  `define AXI_R8_BEA_S16 `i_axi_AXI_R8_BEA_S16
`endif 

`ifdef i_axi_AXI_AR_PYLD_M_W
  `define AXI_AR_PYLD_M_W `i_axi_AXI_AR_PYLD_M_W
`endif 

`ifdef i_axi_AXI_AW_PYLD_M_W
  `define AXI_AW_PYLD_M_W `i_axi_AXI_AW_PYLD_M_W
`endif 

`ifdef i_axi_AXI_W_PYLD_M_W
  `define AXI_W_PYLD_M_W `i_axi_AXI_W_PYLD_M_W
`endif 

`ifdef i_axi_AXI_R_PYLD_M_W
  `define AXI_R_PYLD_M_W `i_axi_AXI_R_PYLD_M_W
`endif 

`ifdef i_axi_AXI_B_PYLD_M_W
  `define AXI_B_PYLD_M_W `i_axi_AXI_B_PYLD_M_W
`endif 

`ifdef i_axi_AXI_AR_PYLD_S_W
  `define AXI_AR_PYLD_S_W `i_axi_AXI_AR_PYLD_S_W
`endif 

`ifdef i_axi_AXI_AW_PYLD_S_W
  `define AXI_AW_PYLD_S_W `i_axi_AXI_AW_PYLD_S_W
`endif 

`ifdef i_axi_AXI_W_PYLD_S_W
  `define AXI_W_PYLD_S_W `i_axi_AXI_W_PYLD_S_W
`endif 

`ifdef i_axi_AXI_R_PYLD_S_W
  `define AXI_R_PYLD_S_W `i_axi_AXI_R_PYLD_S_W
`endif 

`ifdef i_axi_AXI_B_PYLD_S_W
  `define AXI_B_PYLD_S_W `i_axi_AXI_B_PYLD_S_W
`endif 

`ifdef i_axi_AXI_HAS_S0
  `define AXI_HAS_S0 `i_axi_AXI_HAS_S0
`endif 

`ifdef i_axi_AXI_HAS_S1
  `define AXI_HAS_S1 `i_axi_AXI_HAS_S1
`endif 

`ifdef i_axi_AXI_HAS_S2
  `define AXI_HAS_S2 `i_axi_AXI_HAS_S2
`endif 

`ifdef i_axi_AXI_HAS_S3
  `define AXI_HAS_S3 `i_axi_AXI_HAS_S3
`endif 

`ifdef i_axi_AXI_HAS_M1
  `define AXI_HAS_M1 `i_axi_AXI_HAS_M1
`endif 

`ifdef i_axi_AXI_HAS_M2
  `define AXI_HAS_M2 `i_axi_AXI_HAS_M2
`endif 

`ifdef i_axi_AXI_NMV_S0
  `define AXI_NMV_S0 `i_axi_AXI_NMV_S0
`endif 

`ifdef i_axi_AXI_SYS_NUM_FOR_M1
  `define AXI_SYS_NUM_FOR_M1 `i_axi_AXI_SYS_NUM_FOR_M1
`endif 

`ifdef i_axi_AXI_SYS_NUM_FOR_M2
  `define AXI_SYS_NUM_FOR_M2 `i_axi_AXI_SYS_NUM_FOR_M2
`endif 

`ifdef i_axi_AXI_SYS_NUM_FOR_M3
  `define AXI_SYS_NUM_FOR_M3 `i_axi_AXI_SYS_NUM_FOR_M3
`endif 

`ifdef i_axi_AXI_SYS_NUM_FOR_M4
  `define AXI_SYS_NUM_FOR_M4 `i_axi_AXI_SYS_NUM_FOR_M4
`endif 

`ifdef i_axi_AXI_SYS_NUM_FOR_M5
  `define AXI_SYS_NUM_FOR_M5 `i_axi_AXI_SYS_NUM_FOR_M5
`endif 

`ifdef i_axi_AXI_SYS_NUM_FOR_M6
  `define AXI_SYS_NUM_FOR_M6 `i_axi_AXI_SYS_NUM_FOR_M6
`endif 

`ifdef i_axi_AXI_SYS_NUM_FOR_M7
  `define AXI_SYS_NUM_FOR_M7 `i_axi_AXI_SYS_NUM_FOR_M7
`endif 

`ifdef i_axi_AXI_SYS_NUM_FOR_M8
  `define AXI_SYS_NUM_FOR_M8 `i_axi_AXI_SYS_NUM_FOR_M8
`endif 

`ifdef i_axi_AXI_SYS_NUM_FOR_M9
  `define AXI_SYS_NUM_FOR_M9 `i_axi_AXI_SYS_NUM_FOR_M9
`endif 

`ifdef i_axi_AXI_SYS_NUM_FOR_M10
  `define AXI_SYS_NUM_FOR_M10 `i_axi_AXI_SYS_NUM_FOR_M10
`endif 

`ifdef i_axi_AXI_SYS_NUM_FOR_M11
  `define AXI_SYS_NUM_FOR_M11 `i_axi_AXI_SYS_NUM_FOR_M11
`endif 

`ifdef i_axi_AXI_SYS_NUM_FOR_M12
  `define AXI_SYS_NUM_FOR_M12 `i_axi_AXI_SYS_NUM_FOR_M12
`endif 

`ifdef i_axi_AXI_SYS_NUM_FOR_M13
  `define AXI_SYS_NUM_FOR_M13 `i_axi_AXI_SYS_NUM_FOR_M13
`endif 

`ifdef i_axi_AXI_SYS_NUM_FOR_M14
  `define AXI_SYS_NUM_FOR_M14 `i_axi_AXI_SYS_NUM_FOR_M14
`endif 

`ifdef i_axi_AXI_SYS_NUM_FOR_M15
  `define AXI_SYS_NUM_FOR_M15 `i_axi_AXI_SYS_NUM_FOR_M15
`endif 

`ifdef i_axi_AXI_SYS_NUM_FOR_M16
  `define AXI_SYS_NUM_FOR_M16 `i_axi_AXI_SYS_NUM_FOR_M16
`endif 

`ifdef i_axi_AXI_NUM_ICM
  `define AXI_NUM_ICM `i_axi_AXI_NUM_ICM
`endif 

`ifdef i_axi_AXI_ACC_NON_LCL_SLV_S1
  `define AXI_ACC_NON_LCL_SLV_S1 `i_axi_AXI_ACC_NON_LCL_SLV_S1
`endif 

`ifdef i_axi_AXI_ACC_NON_LCL_SLV_S2
  `define AXI_ACC_NON_LCL_SLV_S2 `i_axi_AXI_ACC_NON_LCL_SLV_S2
`endif 

`ifdef i_axi_AXI_ACC_NON_LCL_SLV_S3
  `define AXI_ACC_NON_LCL_SLV_S3 `i_axi_AXI_ACC_NON_LCL_SLV_S3
`endif 

`ifdef i_axi_AXI_ACC_NON_LCL_SLV_S4
  `define AXI_ACC_NON_LCL_SLV_S4 `i_axi_AXI_ACC_NON_LCL_SLV_S4
`endif 

`ifdef i_axi_AXI_ACC_NON_LCL_SLV_S5
  `define AXI_ACC_NON_LCL_SLV_S5 `i_axi_AXI_ACC_NON_LCL_SLV_S5
`endif 

`ifdef i_axi_AXI_ACC_NON_LCL_SLV_S6
  `define AXI_ACC_NON_LCL_SLV_S6 `i_axi_AXI_ACC_NON_LCL_SLV_S6
`endif 

`ifdef i_axi_AXI_ACC_NON_LCL_SLV_S7
  `define AXI_ACC_NON_LCL_SLV_S7 `i_axi_AXI_ACC_NON_LCL_SLV_S7
`endif 

`ifdef i_axi_AXI_ACC_NON_LCL_SLV_S8
  `define AXI_ACC_NON_LCL_SLV_S8 `i_axi_AXI_ACC_NON_LCL_SLV_S8
`endif 

`ifdef i_axi_AXI_ACC_NON_LCL_SLV_S9
  `define AXI_ACC_NON_LCL_SLV_S9 `i_axi_AXI_ACC_NON_LCL_SLV_S9
`endif 

`ifdef i_axi_AXI_ACC_NON_LCL_SLV_S10
  `define AXI_ACC_NON_LCL_SLV_S10 `i_axi_AXI_ACC_NON_LCL_SLV_S10
`endif 

`ifdef i_axi_AXI_ACC_NON_LCL_SLV_S11
  `define AXI_ACC_NON_LCL_SLV_S11 `i_axi_AXI_ACC_NON_LCL_SLV_S11
`endif 

`ifdef i_axi_AXI_ACC_NON_LCL_SLV_S12
  `define AXI_ACC_NON_LCL_SLV_S12 `i_axi_AXI_ACC_NON_LCL_SLV_S12
`endif 

`ifdef i_axi_AXI_ACC_NON_LCL_SLV_S13
  `define AXI_ACC_NON_LCL_SLV_S13 `i_axi_AXI_ACC_NON_LCL_SLV_S13
`endif 

`ifdef i_axi_AXI_ACC_NON_LCL_SLV_S14
  `define AXI_ACC_NON_LCL_SLV_S14 `i_axi_AXI_ACC_NON_LCL_SLV_S14
`endif 

`ifdef i_axi_AXI_ACC_NON_LCL_SLV_S15
  `define AXI_ACC_NON_LCL_SLV_S15 `i_axi_AXI_ACC_NON_LCL_SLV_S15
`endif 

`ifdef i_axi_AXI_ACC_NON_LCL_SLV_S16
  `define AXI_ACC_NON_LCL_SLV_S16 `i_axi_AXI_ACC_NON_LCL_SLV_S16
`endif 

`ifdef i_axi_AXI_IS_ICM_M1
  `define AXI_IS_ICM_M1 `i_axi_AXI_IS_ICM_M1
`endif 

`ifdef i_axi_AXI_IS_ICM_M2
  `define AXI_IS_ICM_M2 `i_axi_AXI_IS_ICM_M2
`endif 

`ifdef i_axi_AXI_IS_ICM_M3
  `define AXI_IS_ICM_M3 `i_axi_AXI_IS_ICM_M3
`endif 

`ifdef i_axi_AXI_IS_ICM_M4
  `define AXI_IS_ICM_M4 `i_axi_AXI_IS_ICM_M4
`endif 

`ifdef i_axi_AXI_IS_ICM_M5
  `define AXI_IS_ICM_M5 `i_axi_AXI_IS_ICM_M5
`endif 

`ifdef i_axi_AXI_IS_ICM_M6
  `define AXI_IS_ICM_M6 `i_axi_AXI_IS_ICM_M6
`endif 

`ifdef i_axi_AXI_IS_ICM_M7
  `define AXI_IS_ICM_M7 `i_axi_AXI_IS_ICM_M7
`endif 

`ifdef i_axi_AXI_IS_ICM_M8
  `define AXI_IS_ICM_M8 `i_axi_AXI_IS_ICM_M8
`endif 

`ifdef i_axi_AXI_IS_ICM_M9
  `define AXI_IS_ICM_M9 `i_axi_AXI_IS_ICM_M9
`endif 

`ifdef i_axi_AXI_IS_ICM_M10
  `define AXI_IS_ICM_M10 `i_axi_AXI_IS_ICM_M10
`endif 

`ifdef i_axi_AXI_IS_ICM_M11
  `define AXI_IS_ICM_M11 `i_axi_AXI_IS_ICM_M11
`endif 

`ifdef i_axi_AXI_IS_ICM_M12
  `define AXI_IS_ICM_M12 `i_axi_AXI_IS_ICM_M12
`endif 

`ifdef i_axi_AXI_IS_ICM_M13
  `define AXI_IS_ICM_M13 `i_axi_AXI_IS_ICM_M13
`endif 

`ifdef i_axi_AXI_IS_ICM_M14
  `define AXI_IS_ICM_M14 `i_axi_AXI_IS_ICM_M14
`endif 

`ifdef i_axi_AXI_IS_ICM_M15
  `define AXI_IS_ICM_M15 `i_axi_AXI_IS_ICM_M15
`endif 

`ifdef i_axi_AXI_IS_ICM_M16
  `define AXI_IS_ICM_M16 `i_axi_AXI_IS_ICM_M16
`endif 

`ifdef i_axi_AXI_HAS_ICM1
  `define AXI_HAS_ICM1 `i_axi_AXI_HAS_ICM1
`endif 

`ifdef i_axi_AXI_HAS_ICM2
  `define AXI_HAS_ICM2 `i_axi_AXI_HAS_ICM2
`endif 

`ifdef i_axi_AXI_HAS_ICM3
  `define AXI_HAS_ICM3 `i_axi_AXI_HAS_ICM3
`endif 

`ifdef i_axi_AXI_HAS_ICM4
  `define AXI_HAS_ICM4 `i_axi_AXI_HAS_ICM4
`endif 

`ifdef i_axi_AXI_IDW_M1
  `define AXI_IDW_M1 `i_axi_AXI_IDW_M1
`endif 

`ifdef i_axi_AXI_IDW_M2
  `define AXI_IDW_M2 `i_axi_AXI_IDW_M2
`endif 

`ifdef i_axi_AXI_IDW_M3
  `define AXI_IDW_M3 `i_axi_AXI_IDW_M3
`endif 

`ifdef i_axi_AXI_IDW_M4
  `define AXI_IDW_M4 `i_axi_AXI_IDW_M4
`endif 

`ifdef i_axi_AXI_NUM_MST_THRU_ICM1
  `define AXI_NUM_MST_THRU_ICM1 `i_axi_AXI_NUM_MST_THRU_ICM1
`endif 

`ifdef i_axi_AXI_NUM_MST_THRU_ICM2
  `define AXI_NUM_MST_THRU_ICM2 `i_axi_AXI_NUM_MST_THRU_ICM2
`endif 

`ifdef i_axi_AXI_NUM_MST_THRU_ICM3
  `define AXI_NUM_MST_THRU_ICM3 `i_axi_AXI_NUM_MST_THRU_ICM3
`endif 

`ifdef i_axi_AXI_NUM_MST_THRU_ICM4
  `define AXI_NUM_MST_THRU_ICM4 `i_axi_AXI_NUM_MST_THRU_ICM4
`endif 

`ifdef i_axi_AXI_ALLOW_MST1_ICM1
  `define AXI_ALLOW_MST1_ICM1 `i_axi_AXI_ALLOW_MST1_ICM1
`endif 

`ifdef i_axi_AXI_ALLOW_MST2_ICM1
  `define AXI_ALLOW_MST2_ICM1 `i_axi_AXI_ALLOW_MST2_ICM1
`endif 

`ifdef i_axi_AXI_ALLOW_MST3_ICM1
  `define AXI_ALLOW_MST3_ICM1 `i_axi_AXI_ALLOW_MST3_ICM1
`endif 

`ifdef i_axi_AXI_ALLOW_MST4_ICM1
  `define AXI_ALLOW_MST4_ICM1 `i_axi_AXI_ALLOW_MST4_ICM1
`endif 

`ifdef i_axi_AXI_ALLOW_MST5_ICM1
  `define AXI_ALLOW_MST5_ICM1 `i_axi_AXI_ALLOW_MST5_ICM1
`endif 

`ifdef i_axi_AXI_ALLOW_MST6_ICM1
  `define AXI_ALLOW_MST6_ICM1 `i_axi_AXI_ALLOW_MST6_ICM1
`endif 

`ifdef i_axi_AXI_ALLOW_MST7_ICM1
  `define AXI_ALLOW_MST7_ICM1 `i_axi_AXI_ALLOW_MST7_ICM1
`endif 

`ifdef i_axi_AXI_ALLOW_MST8_ICM1
  `define AXI_ALLOW_MST8_ICM1 `i_axi_AXI_ALLOW_MST8_ICM1
`endif 

`ifdef i_axi_AXI_ALLOW_MST1_ICM2
  `define AXI_ALLOW_MST1_ICM2 `i_axi_AXI_ALLOW_MST1_ICM2
`endif 

`ifdef i_axi_AXI_ALLOW_MST2_ICM2
  `define AXI_ALLOW_MST2_ICM2 `i_axi_AXI_ALLOW_MST2_ICM2
`endif 

`ifdef i_axi_AXI_ALLOW_MST3_ICM2
  `define AXI_ALLOW_MST3_ICM2 `i_axi_AXI_ALLOW_MST3_ICM2
`endif 

`ifdef i_axi_AXI_ALLOW_MST4_ICM2
  `define AXI_ALLOW_MST4_ICM2 `i_axi_AXI_ALLOW_MST4_ICM2
`endif 

`ifdef i_axi_AXI_ALLOW_MST5_ICM2
  `define AXI_ALLOW_MST5_ICM2 `i_axi_AXI_ALLOW_MST5_ICM2
`endif 

`ifdef i_axi_AXI_ALLOW_MST6_ICM2
  `define AXI_ALLOW_MST6_ICM2 `i_axi_AXI_ALLOW_MST6_ICM2
`endif 

`ifdef i_axi_AXI_ALLOW_MST7_ICM2
  `define AXI_ALLOW_MST7_ICM2 `i_axi_AXI_ALLOW_MST7_ICM2
`endif 

`ifdef i_axi_AXI_ALLOW_MST8_ICM2
  `define AXI_ALLOW_MST8_ICM2 `i_axi_AXI_ALLOW_MST8_ICM2
`endif 

`ifdef i_axi_AXI_ALLOW_MST1_ICM3
  `define AXI_ALLOW_MST1_ICM3 `i_axi_AXI_ALLOW_MST1_ICM3
`endif 

`ifdef i_axi_AXI_ALLOW_MST2_ICM3
  `define AXI_ALLOW_MST2_ICM3 `i_axi_AXI_ALLOW_MST2_ICM3
`endif 

`ifdef i_axi_AXI_ALLOW_MST3_ICM3
  `define AXI_ALLOW_MST3_ICM3 `i_axi_AXI_ALLOW_MST3_ICM3
`endif 

`ifdef i_axi_AXI_ALLOW_MST4_ICM3
  `define AXI_ALLOW_MST4_ICM3 `i_axi_AXI_ALLOW_MST4_ICM3
`endif 

`ifdef i_axi_AXI_ALLOW_MST5_ICM3
  `define AXI_ALLOW_MST5_ICM3 `i_axi_AXI_ALLOW_MST5_ICM3
`endif 

`ifdef i_axi_AXI_ALLOW_MST6_ICM3
  `define AXI_ALLOW_MST6_ICM3 `i_axi_AXI_ALLOW_MST6_ICM3
`endif 

`ifdef i_axi_AXI_ALLOW_MST7_ICM3
  `define AXI_ALLOW_MST7_ICM3 `i_axi_AXI_ALLOW_MST7_ICM3
`endif 

`ifdef i_axi_AXI_ALLOW_MST8_ICM3
  `define AXI_ALLOW_MST8_ICM3 `i_axi_AXI_ALLOW_MST8_ICM3
`endif 

`ifdef i_axi_AXI_ALLOW_MST1_ICM4
  `define AXI_ALLOW_MST1_ICM4 `i_axi_AXI_ALLOW_MST1_ICM4
`endif 

`ifdef i_axi_AXI_ALLOW_MST2_ICM4
  `define AXI_ALLOW_MST2_ICM4 `i_axi_AXI_ALLOW_MST2_ICM4
`endif 

`ifdef i_axi_AXI_ALLOW_MST3_ICM4
  `define AXI_ALLOW_MST3_ICM4 `i_axi_AXI_ALLOW_MST3_ICM4
`endif 

`ifdef i_axi_AXI_ALLOW_MST4_ICM4
  `define AXI_ALLOW_MST4_ICM4 `i_axi_AXI_ALLOW_MST4_ICM4
`endif 

`ifdef i_axi_AXI_ALLOW_MST5_ICM4
  `define AXI_ALLOW_MST5_ICM4 `i_axi_AXI_ALLOW_MST5_ICM4
`endif 

`ifdef i_axi_AXI_ALLOW_MST6_ICM4
  `define AXI_ALLOW_MST6_ICM4 `i_axi_AXI_ALLOW_MST6_ICM4
`endif 

`ifdef i_axi_AXI_ALLOW_MST7_ICM4
  `define AXI_ALLOW_MST7_ICM4 `i_axi_AXI_ALLOW_MST7_ICM4
`endif 

`ifdef i_axi_AXI_ALLOW_MST8_ICM4
  `define AXI_ALLOW_MST8_ICM4 `i_axi_AXI_ALLOW_MST8_ICM4
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M1
  `define AXI_PNUM_FOR_SYS_NUM_M1 `i_axi_AXI_PNUM_FOR_SYS_NUM_M1
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M2
  `define AXI_PNUM_FOR_SYS_NUM_M2 `i_axi_AXI_PNUM_FOR_SYS_NUM_M2
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M3
  `define AXI_PNUM_FOR_SYS_NUM_M3 `i_axi_AXI_PNUM_FOR_SYS_NUM_M3
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M4
  `define AXI_PNUM_FOR_SYS_NUM_M4 `i_axi_AXI_PNUM_FOR_SYS_NUM_M4
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M5
  `define AXI_PNUM_FOR_SYS_NUM_M5 `i_axi_AXI_PNUM_FOR_SYS_NUM_M5
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M6
  `define AXI_PNUM_FOR_SYS_NUM_M6 `i_axi_AXI_PNUM_FOR_SYS_NUM_M6
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M7
  `define AXI_PNUM_FOR_SYS_NUM_M7 `i_axi_AXI_PNUM_FOR_SYS_NUM_M7
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M8
  `define AXI_PNUM_FOR_SYS_NUM_M8 `i_axi_AXI_PNUM_FOR_SYS_NUM_M8
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M9
  `define AXI_PNUM_FOR_SYS_NUM_M9 `i_axi_AXI_PNUM_FOR_SYS_NUM_M9
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M10
  `define AXI_PNUM_FOR_SYS_NUM_M10 `i_axi_AXI_PNUM_FOR_SYS_NUM_M10
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M11
  `define AXI_PNUM_FOR_SYS_NUM_M11 `i_axi_AXI_PNUM_FOR_SYS_NUM_M11
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M12
  `define AXI_PNUM_FOR_SYS_NUM_M12 `i_axi_AXI_PNUM_FOR_SYS_NUM_M12
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M13
  `define AXI_PNUM_FOR_SYS_NUM_M13 `i_axi_AXI_PNUM_FOR_SYS_NUM_M13
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M14
  `define AXI_PNUM_FOR_SYS_NUM_M14 `i_axi_AXI_PNUM_FOR_SYS_NUM_M14
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M15
  `define AXI_PNUM_FOR_SYS_NUM_M15 `i_axi_AXI_PNUM_FOR_SYS_NUM_M15
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M16
  `define AXI_PNUM_FOR_SYS_NUM_M16 `i_axi_AXI_PNUM_FOR_SYS_NUM_M16
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M17
  `define AXI_PNUM_FOR_SYS_NUM_M17 `i_axi_AXI_PNUM_FOR_SYS_NUM_M17
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M18
  `define AXI_PNUM_FOR_SYS_NUM_M18 `i_axi_AXI_PNUM_FOR_SYS_NUM_M18
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M19
  `define AXI_PNUM_FOR_SYS_NUM_M19 `i_axi_AXI_PNUM_FOR_SYS_NUM_M19
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M20
  `define AXI_PNUM_FOR_SYS_NUM_M20 `i_axi_AXI_PNUM_FOR_SYS_NUM_M20
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M21
  `define AXI_PNUM_FOR_SYS_NUM_M21 `i_axi_AXI_PNUM_FOR_SYS_NUM_M21
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M22
  `define AXI_PNUM_FOR_SYS_NUM_M22 `i_axi_AXI_PNUM_FOR_SYS_NUM_M22
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M23
  `define AXI_PNUM_FOR_SYS_NUM_M23 `i_axi_AXI_PNUM_FOR_SYS_NUM_M23
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M24
  `define AXI_PNUM_FOR_SYS_NUM_M24 `i_axi_AXI_PNUM_FOR_SYS_NUM_M24
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M25
  `define AXI_PNUM_FOR_SYS_NUM_M25 `i_axi_AXI_PNUM_FOR_SYS_NUM_M25
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M26
  `define AXI_PNUM_FOR_SYS_NUM_M26 `i_axi_AXI_PNUM_FOR_SYS_NUM_M26
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M27
  `define AXI_PNUM_FOR_SYS_NUM_M27 `i_axi_AXI_PNUM_FOR_SYS_NUM_M27
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M28
  `define AXI_PNUM_FOR_SYS_NUM_M28 `i_axi_AXI_PNUM_FOR_SYS_NUM_M28
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M29
  `define AXI_PNUM_FOR_SYS_NUM_M29 `i_axi_AXI_PNUM_FOR_SYS_NUM_M29
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M30
  `define AXI_PNUM_FOR_SYS_NUM_M30 `i_axi_AXI_PNUM_FOR_SYS_NUM_M30
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M31
  `define AXI_PNUM_FOR_SYS_NUM_M31 `i_axi_AXI_PNUM_FOR_SYS_NUM_M31
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M32
  `define AXI_PNUM_FOR_SYS_NUM_M32 `i_axi_AXI_PNUM_FOR_SYS_NUM_M32
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M33
  `define AXI_PNUM_FOR_SYS_NUM_M33 `i_axi_AXI_PNUM_FOR_SYS_NUM_M33
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M34
  `define AXI_PNUM_FOR_SYS_NUM_M34 `i_axi_AXI_PNUM_FOR_SYS_NUM_M34
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M35
  `define AXI_PNUM_FOR_SYS_NUM_M35 `i_axi_AXI_PNUM_FOR_SYS_NUM_M35
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M36
  `define AXI_PNUM_FOR_SYS_NUM_M36 `i_axi_AXI_PNUM_FOR_SYS_NUM_M36
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M37
  `define AXI_PNUM_FOR_SYS_NUM_M37 `i_axi_AXI_PNUM_FOR_SYS_NUM_M37
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M38
  `define AXI_PNUM_FOR_SYS_NUM_M38 `i_axi_AXI_PNUM_FOR_SYS_NUM_M38
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M39
  `define AXI_PNUM_FOR_SYS_NUM_M39 `i_axi_AXI_PNUM_FOR_SYS_NUM_M39
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M40
  `define AXI_PNUM_FOR_SYS_NUM_M40 `i_axi_AXI_PNUM_FOR_SYS_NUM_M40
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M41
  `define AXI_PNUM_FOR_SYS_NUM_M41 `i_axi_AXI_PNUM_FOR_SYS_NUM_M41
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M42
  `define AXI_PNUM_FOR_SYS_NUM_M42 `i_axi_AXI_PNUM_FOR_SYS_NUM_M42
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M43
  `define AXI_PNUM_FOR_SYS_NUM_M43 `i_axi_AXI_PNUM_FOR_SYS_NUM_M43
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M44
  `define AXI_PNUM_FOR_SYS_NUM_M44 `i_axi_AXI_PNUM_FOR_SYS_NUM_M44
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M45
  `define AXI_PNUM_FOR_SYS_NUM_M45 `i_axi_AXI_PNUM_FOR_SYS_NUM_M45
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M46
  `define AXI_PNUM_FOR_SYS_NUM_M46 `i_axi_AXI_PNUM_FOR_SYS_NUM_M46
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M47
  `define AXI_PNUM_FOR_SYS_NUM_M47 `i_axi_AXI_PNUM_FOR_SYS_NUM_M47
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M48
  `define AXI_PNUM_FOR_SYS_NUM_M48 `i_axi_AXI_PNUM_FOR_SYS_NUM_M48
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M49
  `define AXI_PNUM_FOR_SYS_NUM_M49 `i_axi_AXI_PNUM_FOR_SYS_NUM_M49
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M50
  `define AXI_PNUM_FOR_SYS_NUM_M50 `i_axi_AXI_PNUM_FOR_SYS_NUM_M50
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M51
  `define AXI_PNUM_FOR_SYS_NUM_M51 `i_axi_AXI_PNUM_FOR_SYS_NUM_M51
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M52
  `define AXI_PNUM_FOR_SYS_NUM_M52 `i_axi_AXI_PNUM_FOR_SYS_NUM_M52
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M53
  `define AXI_PNUM_FOR_SYS_NUM_M53 `i_axi_AXI_PNUM_FOR_SYS_NUM_M53
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M54
  `define AXI_PNUM_FOR_SYS_NUM_M54 `i_axi_AXI_PNUM_FOR_SYS_NUM_M54
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M55
  `define AXI_PNUM_FOR_SYS_NUM_M55 `i_axi_AXI_PNUM_FOR_SYS_NUM_M55
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M56
  `define AXI_PNUM_FOR_SYS_NUM_M56 `i_axi_AXI_PNUM_FOR_SYS_NUM_M56
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M57
  `define AXI_PNUM_FOR_SYS_NUM_M57 `i_axi_AXI_PNUM_FOR_SYS_NUM_M57
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M58
  `define AXI_PNUM_FOR_SYS_NUM_M58 `i_axi_AXI_PNUM_FOR_SYS_NUM_M58
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M59
  `define AXI_PNUM_FOR_SYS_NUM_M59 `i_axi_AXI_PNUM_FOR_SYS_NUM_M59
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M60
  `define AXI_PNUM_FOR_SYS_NUM_M60 `i_axi_AXI_PNUM_FOR_SYS_NUM_M60
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M61
  `define AXI_PNUM_FOR_SYS_NUM_M61 `i_axi_AXI_PNUM_FOR_SYS_NUM_M61
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M62
  `define AXI_PNUM_FOR_SYS_NUM_M62 `i_axi_AXI_PNUM_FOR_SYS_NUM_M62
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M63
  `define AXI_PNUM_FOR_SYS_NUM_M63 `i_axi_AXI_PNUM_FOR_SYS_NUM_M63
`endif 

`ifdef i_axi_AXI_PNUM_FOR_SYS_NUM_M64
  `define AXI_PNUM_FOR_SYS_NUM_M64 `i_axi_AXI_PNUM_FOR_SYS_NUM_M64
`endif 

`ifdef i_axi_AXI_QOS
  `define AXI_QOS `i_axi_AXI_QOS
`endif 

`ifdef i_axi_AXI_SRC_LICENSE_CHK
  `define AXI_SRC_LICENSE_CHK `i_axi_AXI_SRC_LICENSE_CHK
`endif 

`ifdef i_axi_AXI_NSPV_M1_AR_QOSARB
  `define AXI_NSPV_M1_AR_QOSARB `i_axi_AXI_NSPV_M1_AR_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M2_AR_QOSARB
  `define AXI_NSPV_M2_AR_QOSARB `i_axi_AXI_NSPV_M2_AR_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M3_AR_QOSARB
  `define AXI_NSPV_M3_AR_QOSARB `i_axi_AXI_NSPV_M3_AR_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M4_AR_QOSARB
  `define AXI_NSPV_M4_AR_QOSARB `i_axi_AXI_NSPV_M4_AR_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M5_AR_QOSARB
  `define AXI_NSPV_M5_AR_QOSARB `i_axi_AXI_NSPV_M5_AR_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M6_AR_QOSARB
  `define AXI_NSPV_M6_AR_QOSARB `i_axi_AXI_NSPV_M6_AR_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M7_AR_QOSARB
  `define AXI_NSPV_M7_AR_QOSARB `i_axi_AXI_NSPV_M7_AR_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M8_AR_QOSARB
  `define AXI_NSPV_M8_AR_QOSARB `i_axi_AXI_NSPV_M8_AR_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M9_AR_QOSARB
  `define AXI_NSPV_M9_AR_QOSARB `i_axi_AXI_NSPV_M9_AR_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M10_AR_QOSARB
  `define AXI_NSPV_M10_AR_QOSARB `i_axi_AXI_NSPV_M10_AR_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M11_AR_QOSARB
  `define AXI_NSPV_M11_AR_QOSARB `i_axi_AXI_NSPV_M11_AR_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M12_AR_QOSARB
  `define AXI_NSPV_M12_AR_QOSARB `i_axi_AXI_NSPV_M12_AR_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M13_AR_QOSARB
  `define AXI_NSPV_M13_AR_QOSARB `i_axi_AXI_NSPV_M13_AR_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M14_AR_QOSARB
  `define AXI_NSPV_M14_AR_QOSARB `i_axi_AXI_NSPV_M14_AR_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M15_AR_QOSARB
  `define AXI_NSPV_M15_AR_QOSARB `i_axi_AXI_NSPV_M15_AR_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M16_AR_QOSARB
  `define AXI_NSPV_M16_AR_QOSARB `i_axi_AXI_NSPV_M16_AR_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M1_AW_QOSARB
  `define AXI_NSPV_M1_AW_QOSARB `i_axi_AXI_NSPV_M1_AW_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M2_AW_QOSARB
  `define AXI_NSPV_M2_AW_QOSARB `i_axi_AXI_NSPV_M2_AW_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M3_AW_QOSARB
  `define AXI_NSPV_M3_AW_QOSARB `i_axi_AXI_NSPV_M3_AW_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M4_AW_QOSARB
  `define AXI_NSPV_M4_AW_QOSARB `i_axi_AXI_NSPV_M4_AW_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M5_AW_QOSARB
  `define AXI_NSPV_M5_AW_QOSARB `i_axi_AXI_NSPV_M5_AW_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M6_AW_QOSARB
  `define AXI_NSPV_M6_AW_QOSARB `i_axi_AXI_NSPV_M6_AW_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M7_AW_QOSARB
  `define AXI_NSPV_M7_AW_QOSARB `i_axi_AXI_NSPV_M7_AW_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M8_AW_QOSARB
  `define AXI_NSPV_M8_AW_QOSARB `i_axi_AXI_NSPV_M8_AW_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M9_AW_QOSARB
  `define AXI_NSPV_M9_AW_QOSARB `i_axi_AXI_NSPV_M9_AW_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M10_AW_QOSARB
  `define AXI_NSPV_M10_AW_QOSARB `i_axi_AXI_NSPV_M10_AW_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M11_AW_QOSARB
  `define AXI_NSPV_M11_AW_QOSARB `i_axi_AXI_NSPV_M11_AW_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M12_AW_QOSARB
  `define AXI_NSPV_M12_AW_QOSARB `i_axi_AXI_NSPV_M12_AW_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M13_AW_QOSARB
  `define AXI_NSPV_M13_AW_QOSARB `i_axi_AXI_NSPV_M13_AW_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M14_AW_QOSARB
  `define AXI_NSPV_M14_AW_QOSARB `i_axi_AXI_NSPV_M14_AW_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M15_AW_QOSARB
  `define AXI_NSPV_M15_AW_QOSARB `i_axi_AXI_NSPV_M15_AW_QOSARB
`endif 

`ifdef i_axi_AXI_NSPV_M16_AW_QOSARB
  `define AXI_NSPV_M16_AW_QOSARB `i_axi_AXI_NSPV_M16_AW_QOSARB
`endif 

`ifdef i_axi_AXI_AR_HAS_QOS_REGULATOR_M1
  `define AXI_AR_HAS_QOS_REGULATOR_M1 `i_axi_AXI_AR_HAS_QOS_REGULATOR_M1
`endif 

`ifdef i_axi_AXI_AR_QOS_REGULATOR_M1
  `define AXI_AR_QOS_REGULATOR_M1 `i_axi_AXI_AR_QOS_REGULATOR_M1
`endif 

`ifdef i_axi_AXI_AR_HAS_QOS_REGULATOR_M2
  `define AXI_AR_HAS_QOS_REGULATOR_M2 `i_axi_AXI_AR_HAS_QOS_REGULATOR_M2
`endif 

`ifdef i_axi_AXI_AR_QOS_REGULATOR_M2
  `define AXI_AR_QOS_REGULATOR_M2 `i_axi_AXI_AR_QOS_REGULATOR_M2
`endif 

`ifdef i_axi_AXI_AR_HAS_QOS_REGULATOR_M3
  `define AXI_AR_HAS_QOS_REGULATOR_M3 `i_axi_AXI_AR_HAS_QOS_REGULATOR_M3
`endif 

`ifdef i_axi_AXI_AR_QOS_REGULATOR_M3
  `define AXI_AR_QOS_REGULATOR_M3 `i_axi_AXI_AR_QOS_REGULATOR_M3
`endif 

`ifdef i_axi_AXI_AR_HAS_QOS_REGULATOR_M4
  `define AXI_AR_HAS_QOS_REGULATOR_M4 `i_axi_AXI_AR_HAS_QOS_REGULATOR_M4
`endif 

`ifdef i_axi_AXI_AR_QOS_REGULATOR_M4
  `define AXI_AR_QOS_REGULATOR_M4 `i_axi_AXI_AR_QOS_REGULATOR_M4
`endif 

`ifdef i_axi_AXI_AR_HAS_QOS_REGULATOR_M5
  `define AXI_AR_HAS_QOS_REGULATOR_M5 `i_axi_AXI_AR_HAS_QOS_REGULATOR_M5
`endif 

`ifdef i_axi_AXI_AR_QOS_REGULATOR_M5
  `define AXI_AR_QOS_REGULATOR_M5 `i_axi_AXI_AR_QOS_REGULATOR_M5
`endif 

`ifdef i_axi_AXI_AR_HAS_QOS_REGULATOR_M6
  `define AXI_AR_HAS_QOS_REGULATOR_M6 `i_axi_AXI_AR_HAS_QOS_REGULATOR_M6
`endif 

`ifdef i_axi_AXI_AR_QOS_REGULATOR_M6
  `define AXI_AR_QOS_REGULATOR_M6 `i_axi_AXI_AR_QOS_REGULATOR_M6
`endif 

`ifdef i_axi_AXI_AR_HAS_QOS_REGULATOR_M7
  `define AXI_AR_HAS_QOS_REGULATOR_M7 `i_axi_AXI_AR_HAS_QOS_REGULATOR_M7
`endif 

`ifdef i_axi_AXI_AR_QOS_REGULATOR_M7
  `define AXI_AR_QOS_REGULATOR_M7 `i_axi_AXI_AR_QOS_REGULATOR_M7
`endif 

`ifdef i_axi_AXI_AR_HAS_QOS_REGULATOR_M8
  `define AXI_AR_HAS_QOS_REGULATOR_M8 `i_axi_AXI_AR_HAS_QOS_REGULATOR_M8
`endif 

`ifdef i_axi_AXI_AR_QOS_REGULATOR_M8
  `define AXI_AR_QOS_REGULATOR_M8 `i_axi_AXI_AR_QOS_REGULATOR_M8
`endif 

`ifdef i_axi_AXI_AR_HAS_QOS_REGULATOR_M9
  `define AXI_AR_HAS_QOS_REGULATOR_M9 `i_axi_AXI_AR_HAS_QOS_REGULATOR_M9
`endif 

`ifdef i_axi_AXI_AR_QOS_REGULATOR_M9
  `define AXI_AR_QOS_REGULATOR_M9 `i_axi_AXI_AR_QOS_REGULATOR_M9
`endif 

`ifdef i_axi_AXI_AR_HAS_QOS_REGULATOR_M10
  `define AXI_AR_HAS_QOS_REGULATOR_M10 `i_axi_AXI_AR_HAS_QOS_REGULATOR_M10
`endif 

`ifdef i_axi_AXI_AR_QOS_REGULATOR_M10
  `define AXI_AR_QOS_REGULATOR_M10 `i_axi_AXI_AR_QOS_REGULATOR_M10
`endif 

`ifdef i_axi_AXI_AR_HAS_QOS_REGULATOR_M11
  `define AXI_AR_HAS_QOS_REGULATOR_M11 `i_axi_AXI_AR_HAS_QOS_REGULATOR_M11
`endif 

`ifdef i_axi_AXI_AR_QOS_REGULATOR_M11
  `define AXI_AR_QOS_REGULATOR_M11 `i_axi_AXI_AR_QOS_REGULATOR_M11
`endif 

`ifdef i_axi_AXI_AR_HAS_QOS_REGULATOR_M12
  `define AXI_AR_HAS_QOS_REGULATOR_M12 `i_axi_AXI_AR_HAS_QOS_REGULATOR_M12
`endif 

`ifdef i_axi_AXI_AR_QOS_REGULATOR_M12
  `define AXI_AR_QOS_REGULATOR_M12 `i_axi_AXI_AR_QOS_REGULATOR_M12
`endif 

`ifdef i_axi_AXI_AR_HAS_QOS_REGULATOR_M13
  `define AXI_AR_HAS_QOS_REGULATOR_M13 `i_axi_AXI_AR_HAS_QOS_REGULATOR_M13
`endif 

`ifdef i_axi_AXI_AR_QOS_REGULATOR_M13
  `define AXI_AR_QOS_REGULATOR_M13 `i_axi_AXI_AR_QOS_REGULATOR_M13
`endif 

`ifdef i_axi_AXI_AR_HAS_QOS_REGULATOR_M14
  `define AXI_AR_HAS_QOS_REGULATOR_M14 `i_axi_AXI_AR_HAS_QOS_REGULATOR_M14
`endif 

`ifdef i_axi_AXI_AR_QOS_REGULATOR_M14
  `define AXI_AR_QOS_REGULATOR_M14 `i_axi_AXI_AR_QOS_REGULATOR_M14
`endif 

`ifdef i_axi_AXI_AR_HAS_QOS_REGULATOR_M15
  `define AXI_AR_HAS_QOS_REGULATOR_M15 `i_axi_AXI_AR_HAS_QOS_REGULATOR_M15
`endif 

`ifdef i_axi_AXI_AR_QOS_REGULATOR_M15
  `define AXI_AR_QOS_REGULATOR_M15 `i_axi_AXI_AR_QOS_REGULATOR_M15
`endif 

`ifdef i_axi_AXI_AR_HAS_QOS_REGULATOR_M16
  `define AXI_AR_HAS_QOS_REGULATOR_M16 `i_axi_AXI_AR_HAS_QOS_REGULATOR_M16
`endif 

`ifdef i_axi_AXI_AR_QOS_REGULATOR_M16
  `define AXI_AR_QOS_REGULATOR_M16 `i_axi_AXI_AR_QOS_REGULATOR_M16
`endif 

`ifdef i_axi_AXI_AW_HAS_QOS_REGULATOR_M1
  `define AXI_AW_HAS_QOS_REGULATOR_M1 `i_axi_AXI_AW_HAS_QOS_REGULATOR_M1
`endif 

`ifdef i_axi_AXI_AW_QOS_REGULATOR_M1
  `define AXI_AW_QOS_REGULATOR_M1 `i_axi_AXI_AW_QOS_REGULATOR_M1
`endif 

`ifdef i_axi_AXI_AW_HAS_QOS_REGULATOR_M2
  `define AXI_AW_HAS_QOS_REGULATOR_M2 `i_axi_AXI_AW_HAS_QOS_REGULATOR_M2
`endif 

`ifdef i_axi_AXI_AW_QOS_REGULATOR_M2
  `define AXI_AW_QOS_REGULATOR_M2 `i_axi_AXI_AW_QOS_REGULATOR_M2
`endif 

`ifdef i_axi_AXI_AW_HAS_QOS_REGULATOR_M3
  `define AXI_AW_HAS_QOS_REGULATOR_M3 `i_axi_AXI_AW_HAS_QOS_REGULATOR_M3
`endif 

`ifdef i_axi_AXI_AW_QOS_REGULATOR_M3
  `define AXI_AW_QOS_REGULATOR_M3 `i_axi_AXI_AW_QOS_REGULATOR_M3
`endif 

`ifdef i_axi_AXI_AW_HAS_QOS_REGULATOR_M4
  `define AXI_AW_HAS_QOS_REGULATOR_M4 `i_axi_AXI_AW_HAS_QOS_REGULATOR_M4
`endif 

`ifdef i_axi_AXI_AW_QOS_REGULATOR_M4
  `define AXI_AW_QOS_REGULATOR_M4 `i_axi_AXI_AW_QOS_REGULATOR_M4
`endif 

`ifdef i_axi_AXI_AW_HAS_QOS_REGULATOR_M5
  `define AXI_AW_HAS_QOS_REGULATOR_M5 `i_axi_AXI_AW_HAS_QOS_REGULATOR_M5
`endif 

`ifdef i_axi_AXI_AW_QOS_REGULATOR_M5
  `define AXI_AW_QOS_REGULATOR_M5 `i_axi_AXI_AW_QOS_REGULATOR_M5
`endif 

`ifdef i_axi_AXI_AW_HAS_QOS_REGULATOR_M6
  `define AXI_AW_HAS_QOS_REGULATOR_M6 `i_axi_AXI_AW_HAS_QOS_REGULATOR_M6
`endif 

`ifdef i_axi_AXI_AW_QOS_REGULATOR_M6
  `define AXI_AW_QOS_REGULATOR_M6 `i_axi_AXI_AW_QOS_REGULATOR_M6
`endif 

`ifdef i_axi_AXI_AW_HAS_QOS_REGULATOR_M7
  `define AXI_AW_HAS_QOS_REGULATOR_M7 `i_axi_AXI_AW_HAS_QOS_REGULATOR_M7
`endif 

`ifdef i_axi_AXI_AW_QOS_REGULATOR_M7
  `define AXI_AW_QOS_REGULATOR_M7 `i_axi_AXI_AW_QOS_REGULATOR_M7
`endif 

`ifdef i_axi_AXI_AW_HAS_QOS_REGULATOR_M8
  `define AXI_AW_HAS_QOS_REGULATOR_M8 `i_axi_AXI_AW_HAS_QOS_REGULATOR_M8
`endif 

`ifdef i_axi_AXI_AW_QOS_REGULATOR_M8
  `define AXI_AW_QOS_REGULATOR_M8 `i_axi_AXI_AW_QOS_REGULATOR_M8
`endif 

`ifdef i_axi_AXI_AW_HAS_QOS_REGULATOR_M9
  `define AXI_AW_HAS_QOS_REGULATOR_M9 `i_axi_AXI_AW_HAS_QOS_REGULATOR_M9
`endif 

`ifdef i_axi_AXI_AW_QOS_REGULATOR_M9
  `define AXI_AW_QOS_REGULATOR_M9 `i_axi_AXI_AW_QOS_REGULATOR_M9
`endif 

`ifdef i_axi_AXI_AW_HAS_QOS_REGULATOR_M10
  `define AXI_AW_HAS_QOS_REGULATOR_M10 `i_axi_AXI_AW_HAS_QOS_REGULATOR_M10
`endif 

`ifdef i_axi_AXI_AW_QOS_REGULATOR_M10
  `define AXI_AW_QOS_REGULATOR_M10 `i_axi_AXI_AW_QOS_REGULATOR_M10
`endif 

`ifdef i_axi_AXI_AW_HAS_QOS_REGULATOR_M11
  `define AXI_AW_HAS_QOS_REGULATOR_M11 `i_axi_AXI_AW_HAS_QOS_REGULATOR_M11
`endif 

`ifdef i_axi_AXI_AW_QOS_REGULATOR_M11
  `define AXI_AW_QOS_REGULATOR_M11 `i_axi_AXI_AW_QOS_REGULATOR_M11
`endif 

`ifdef i_axi_AXI_AW_HAS_QOS_REGULATOR_M12
  `define AXI_AW_HAS_QOS_REGULATOR_M12 `i_axi_AXI_AW_HAS_QOS_REGULATOR_M12
`endif 

`ifdef i_axi_AXI_AW_QOS_REGULATOR_M12
  `define AXI_AW_QOS_REGULATOR_M12 `i_axi_AXI_AW_QOS_REGULATOR_M12
`endif 

`ifdef i_axi_AXI_AW_HAS_QOS_REGULATOR_M13
  `define AXI_AW_HAS_QOS_REGULATOR_M13 `i_axi_AXI_AW_HAS_QOS_REGULATOR_M13
`endif 

`ifdef i_axi_AXI_AW_QOS_REGULATOR_M13
  `define AXI_AW_QOS_REGULATOR_M13 `i_axi_AXI_AW_QOS_REGULATOR_M13
`endif 

`ifdef i_axi_AXI_AW_HAS_QOS_REGULATOR_M14
  `define AXI_AW_HAS_QOS_REGULATOR_M14 `i_axi_AXI_AW_HAS_QOS_REGULATOR_M14
`endif 

`ifdef i_axi_AXI_AW_QOS_REGULATOR_M14
  `define AXI_AW_QOS_REGULATOR_M14 `i_axi_AXI_AW_QOS_REGULATOR_M14
`endif 

`ifdef i_axi_AXI_AW_HAS_QOS_REGULATOR_M15
  `define AXI_AW_HAS_QOS_REGULATOR_M15 `i_axi_AXI_AW_HAS_QOS_REGULATOR_M15
`endif 

`ifdef i_axi_AXI_AW_QOS_REGULATOR_M15
  `define AXI_AW_QOS_REGULATOR_M15 `i_axi_AXI_AW_QOS_REGULATOR_M15
`endif 

`ifdef i_axi_AXI_AW_HAS_QOS_REGULATOR_M16
  `define AXI_AW_HAS_QOS_REGULATOR_M16 `i_axi_AXI_AW_HAS_QOS_REGULATOR_M16
`endif 

`ifdef i_axi_AXI_AW_QOS_REGULATOR_M16
  `define AXI_AW_QOS_REGULATOR_M16 `i_axi_AXI_AW_QOS_REGULATOR_M16
`endif 

`ifdef i_axi_AXI_HAS_ARQOS_EXT_M1
  `define AXI_HAS_ARQOS_EXT_M1 `i_axi_AXI_HAS_ARQOS_EXT_M1
`endif 

`ifdef i_axi_AXI_ARQOS_EXT_M1
  `define AXI_ARQOS_EXT_M1 `i_axi_AXI_ARQOS_EXT_M1
`endif 

`ifdef i_axi_AXI_ARQOS_INT_M1
  `define AXI_ARQOS_INT_M1 `i_axi_AXI_ARQOS_INT_M1
`endif 

`ifdef i_axi_AXI_HAS_ARQOS_EXT_M2
  `define AXI_HAS_ARQOS_EXT_M2 `i_axi_AXI_HAS_ARQOS_EXT_M2
`endif 

`ifdef i_axi_AXI_ARQOS_EXT_M2
  `define AXI_ARQOS_EXT_M2 `i_axi_AXI_ARQOS_EXT_M2
`endif 

`ifdef i_axi_AXI_ARQOS_INT_M2
  `define AXI_ARQOS_INT_M2 `i_axi_AXI_ARQOS_INT_M2
`endif 

`ifdef i_axi_AXI_HAS_ARQOS_EXT_M3
  `define AXI_HAS_ARQOS_EXT_M3 `i_axi_AXI_HAS_ARQOS_EXT_M3
`endif 

`ifdef i_axi_AXI_ARQOS_EXT_M3
  `define AXI_ARQOS_EXT_M3 `i_axi_AXI_ARQOS_EXT_M3
`endif 

`ifdef i_axi_AXI_ARQOS_INT_M3
  `define AXI_ARQOS_INT_M3 `i_axi_AXI_ARQOS_INT_M3
`endif 

`ifdef i_axi_AXI_HAS_ARQOS_EXT_M4
  `define AXI_HAS_ARQOS_EXT_M4 `i_axi_AXI_HAS_ARQOS_EXT_M4
`endif 

`ifdef i_axi_AXI_ARQOS_EXT_M4
  `define AXI_ARQOS_EXT_M4 `i_axi_AXI_ARQOS_EXT_M4
`endif 

`ifdef i_axi_AXI_ARQOS_INT_M4
  `define AXI_ARQOS_INT_M4 `i_axi_AXI_ARQOS_INT_M4
`endif 

`ifdef i_axi_AXI_HAS_ARQOS_EXT_M5
  `define AXI_HAS_ARQOS_EXT_M5 `i_axi_AXI_HAS_ARQOS_EXT_M5
`endif 

`ifdef i_axi_AXI_ARQOS_EXT_M5
  `define AXI_ARQOS_EXT_M5 `i_axi_AXI_ARQOS_EXT_M5
`endif 

`ifdef i_axi_AXI_ARQOS_INT_M5
  `define AXI_ARQOS_INT_M5 `i_axi_AXI_ARQOS_INT_M5
`endif 

`ifdef i_axi_AXI_HAS_ARQOS_EXT_M6
  `define AXI_HAS_ARQOS_EXT_M6 `i_axi_AXI_HAS_ARQOS_EXT_M6
`endif 

`ifdef i_axi_AXI_ARQOS_EXT_M6
  `define AXI_ARQOS_EXT_M6 `i_axi_AXI_ARQOS_EXT_M6
`endif 

`ifdef i_axi_AXI_ARQOS_INT_M6
  `define AXI_ARQOS_INT_M6 `i_axi_AXI_ARQOS_INT_M6
`endif 

`ifdef i_axi_AXI_HAS_ARQOS_EXT_M7
  `define AXI_HAS_ARQOS_EXT_M7 `i_axi_AXI_HAS_ARQOS_EXT_M7
`endif 

`ifdef i_axi_AXI_ARQOS_EXT_M7
  `define AXI_ARQOS_EXT_M7 `i_axi_AXI_ARQOS_EXT_M7
`endif 

`ifdef i_axi_AXI_ARQOS_INT_M7
  `define AXI_ARQOS_INT_M7 `i_axi_AXI_ARQOS_INT_M7
`endif 

`ifdef i_axi_AXI_HAS_ARQOS_EXT_M8
  `define AXI_HAS_ARQOS_EXT_M8 `i_axi_AXI_HAS_ARQOS_EXT_M8
`endif 

`ifdef i_axi_AXI_ARQOS_EXT_M8
  `define AXI_ARQOS_EXT_M8 `i_axi_AXI_ARQOS_EXT_M8
`endif 

`ifdef i_axi_AXI_ARQOS_INT_M8
  `define AXI_ARQOS_INT_M8 `i_axi_AXI_ARQOS_INT_M8
`endif 

`ifdef i_axi_AXI_HAS_ARQOS_EXT_M9
  `define AXI_HAS_ARQOS_EXT_M9 `i_axi_AXI_HAS_ARQOS_EXT_M9
`endif 

`ifdef i_axi_AXI_ARQOS_EXT_M9
  `define AXI_ARQOS_EXT_M9 `i_axi_AXI_ARQOS_EXT_M9
`endif 

`ifdef i_axi_AXI_ARQOS_INT_M9
  `define AXI_ARQOS_INT_M9 `i_axi_AXI_ARQOS_INT_M9
`endif 

`ifdef i_axi_AXI_HAS_ARQOS_EXT_M10
  `define AXI_HAS_ARQOS_EXT_M10 `i_axi_AXI_HAS_ARQOS_EXT_M10
`endif 

`ifdef i_axi_AXI_ARQOS_EXT_M10
  `define AXI_ARQOS_EXT_M10 `i_axi_AXI_ARQOS_EXT_M10
`endif 

`ifdef i_axi_AXI_ARQOS_INT_M10
  `define AXI_ARQOS_INT_M10 `i_axi_AXI_ARQOS_INT_M10
`endif 

`ifdef i_axi_AXI_HAS_ARQOS_EXT_M11
  `define AXI_HAS_ARQOS_EXT_M11 `i_axi_AXI_HAS_ARQOS_EXT_M11
`endif 

`ifdef i_axi_AXI_ARQOS_EXT_M11
  `define AXI_ARQOS_EXT_M11 `i_axi_AXI_ARQOS_EXT_M11
`endif 

`ifdef i_axi_AXI_ARQOS_INT_M11
  `define AXI_ARQOS_INT_M11 `i_axi_AXI_ARQOS_INT_M11
`endif 

`ifdef i_axi_AXI_HAS_ARQOS_EXT_M12
  `define AXI_HAS_ARQOS_EXT_M12 `i_axi_AXI_HAS_ARQOS_EXT_M12
`endif 

`ifdef i_axi_AXI_ARQOS_EXT_M12
  `define AXI_ARQOS_EXT_M12 `i_axi_AXI_ARQOS_EXT_M12
`endif 

`ifdef i_axi_AXI_ARQOS_INT_M12
  `define AXI_ARQOS_INT_M12 `i_axi_AXI_ARQOS_INT_M12
`endif 

`ifdef i_axi_AXI_HAS_ARQOS_EXT_M13
  `define AXI_HAS_ARQOS_EXT_M13 `i_axi_AXI_HAS_ARQOS_EXT_M13
`endif 

`ifdef i_axi_AXI_ARQOS_EXT_M13
  `define AXI_ARQOS_EXT_M13 `i_axi_AXI_ARQOS_EXT_M13
`endif 

`ifdef i_axi_AXI_ARQOS_INT_M13
  `define AXI_ARQOS_INT_M13 `i_axi_AXI_ARQOS_INT_M13
`endif 

`ifdef i_axi_AXI_HAS_ARQOS_EXT_M14
  `define AXI_HAS_ARQOS_EXT_M14 `i_axi_AXI_HAS_ARQOS_EXT_M14
`endif 

`ifdef i_axi_AXI_ARQOS_EXT_M14
  `define AXI_ARQOS_EXT_M14 `i_axi_AXI_ARQOS_EXT_M14
`endif 

`ifdef i_axi_AXI_ARQOS_INT_M14
  `define AXI_ARQOS_INT_M14 `i_axi_AXI_ARQOS_INT_M14
`endif 

`ifdef i_axi_AXI_HAS_ARQOS_EXT_M15
  `define AXI_HAS_ARQOS_EXT_M15 `i_axi_AXI_HAS_ARQOS_EXT_M15
`endif 

`ifdef i_axi_AXI_ARQOS_EXT_M15
  `define AXI_ARQOS_EXT_M15 `i_axi_AXI_ARQOS_EXT_M15
`endif 

`ifdef i_axi_AXI_ARQOS_INT_M15
  `define AXI_ARQOS_INT_M15 `i_axi_AXI_ARQOS_INT_M15
`endif 

`ifdef i_axi_AXI_HAS_ARQOS_EXT_M16
  `define AXI_HAS_ARQOS_EXT_M16 `i_axi_AXI_HAS_ARQOS_EXT_M16
`endif 

`ifdef i_axi_AXI_ARQOS_EXT_M16
  `define AXI_ARQOS_EXT_M16 `i_axi_AXI_ARQOS_EXT_M16
`endif 

`ifdef i_axi_AXI_ARQOS_INT_M16
  `define AXI_ARQOS_INT_M16 `i_axi_AXI_ARQOS_INT_M16
`endif 

`ifdef i_axi_AXI_HAS_AWQOS_EXT_M1
  `define AXI_HAS_AWQOS_EXT_M1 `i_axi_AXI_HAS_AWQOS_EXT_M1
`endif 

`ifdef i_axi_AXI_AWQOS_EXT_M1
  `define AXI_AWQOS_EXT_M1 `i_axi_AXI_AWQOS_EXT_M1
`endif 

`ifdef i_axi_AXI_AWQOS_INT_M1
  `define AXI_AWQOS_INT_M1 `i_axi_AXI_AWQOS_INT_M1
`endif 

`ifdef i_axi_AXI_HAS_AWQOS_EXT_M2
  `define AXI_HAS_AWQOS_EXT_M2 `i_axi_AXI_HAS_AWQOS_EXT_M2
`endif 

`ifdef i_axi_AXI_AWQOS_EXT_M2
  `define AXI_AWQOS_EXT_M2 `i_axi_AXI_AWQOS_EXT_M2
`endif 

`ifdef i_axi_AXI_AWQOS_INT_M2
  `define AXI_AWQOS_INT_M2 `i_axi_AXI_AWQOS_INT_M2
`endif 

`ifdef i_axi_AXI_HAS_AWQOS_EXT_M3
  `define AXI_HAS_AWQOS_EXT_M3 `i_axi_AXI_HAS_AWQOS_EXT_M3
`endif 

`ifdef i_axi_AXI_AWQOS_EXT_M3
  `define AXI_AWQOS_EXT_M3 `i_axi_AXI_AWQOS_EXT_M3
`endif 

`ifdef i_axi_AXI_AWQOS_INT_M3
  `define AXI_AWQOS_INT_M3 `i_axi_AXI_AWQOS_INT_M3
`endif 

`ifdef i_axi_AXI_HAS_AWQOS_EXT_M4
  `define AXI_HAS_AWQOS_EXT_M4 `i_axi_AXI_HAS_AWQOS_EXT_M4
`endif 

`ifdef i_axi_AXI_AWQOS_EXT_M4
  `define AXI_AWQOS_EXT_M4 `i_axi_AXI_AWQOS_EXT_M4
`endif 

`ifdef i_axi_AXI_AWQOS_INT_M4
  `define AXI_AWQOS_INT_M4 `i_axi_AXI_AWQOS_INT_M4
`endif 

`ifdef i_axi_AXI_HAS_AWQOS_EXT_M5
  `define AXI_HAS_AWQOS_EXT_M5 `i_axi_AXI_HAS_AWQOS_EXT_M5
`endif 

`ifdef i_axi_AXI_AWQOS_EXT_M5
  `define AXI_AWQOS_EXT_M5 `i_axi_AXI_AWQOS_EXT_M5
`endif 

`ifdef i_axi_AXI_AWQOS_INT_M5
  `define AXI_AWQOS_INT_M5 `i_axi_AXI_AWQOS_INT_M5
`endif 

`ifdef i_axi_AXI_HAS_AWQOS_EXT_M6
  `define AXI_HAS_AWQOS_EXT_M6 `i_axi_AXI_HAS_AWQOS_EXT_M6
`endif 

`ifdef i_axi_AXI_AWQOS_EXT_M6
  `define AXI_AWQOS_EXT_M6 `i_axi_AXI_AWQOS_EXT_M6
`endif 

`ifdef i_axi_AXI_AWQOS_INT_M6
  `define AXI_AWQOS_INT_M6 `i_axi_AXI_AWQOS_INT_M6
`endif 

`ifdef i_axi_AXI_HAS_AWQOS_EXT_M7
  `define AXI_HAS_AWQOS_EXT_M7 `i_axi_AXI_HAS_AWQOS_EXT_M7
`endif 

`ifdef i_axi_AXI_AWQOS_EXT_M7
  `define AXI_AWQOS_EXT_M7 `i_axi_AXI_AWQOS_EXT_M7
`endif 

`ifdef i_axi_AXI_AWQOS_INT_M7
  `define AXI_AWQOS_INT_M7 `i_axi_AXI_AWQOS_INT_M7
`endif 

`ifdef i_axi_AXI_HAS_AWQOS_EXT_M8
  `define AXI_HAS_AWQOS_EXT_M8 `i_axi_AXI_HAS_AWQOS_EXT_M8
`endif 

`ifdef i_axi_AXI_AWQOS_EXT_M8
  `define AXI_AWQOS_EXT_M8 `i_axi_AXI_AWQOS_EXT_M8
`endif 

`ifdef i_axi_AXI_AWQOS_INT_M8
  `define AXI_AWQOS_INT_M8 `i_axi_AXI_AWQOS_INT_M8
`endif 

`ifdef i_axi_AXI_HAS_AWQOS_EXT_M9
  `define AXI_HAS_AWQOS_EXT_M9 `i_axi_AXI_HAS_AWQOS_EXT_M9
`endif 

`ifdef i_axi_AXI_AWQOS_EXT_M9
  `define AXI_AWQOS_EXT_M9 `i_axi_AXI_AWQOS_EXT_M9
`endif 

`ifdef i_axi_AXI_AWQOS_INT_M9
  `define AXI_AWQOS_INT_M9 `i_axi_AXI_AWQOS_INT_M9
`endif 

`ifdef i_axi_AXI_HAS_AWQOS_EXT_M10
  `define AXI_HAS_AWQOS_EXT_M10 `i_axi_AXI_HAS_AWQOS_EXT_M10
`endif 

`ifdef i_axi_AXI_AWQOS_EXT_M10
  `define AXI_AWQOS_EXT_M10 `i_axi_AXI_AWQOS_EXT_M10
`endif 

`ifdef i_axi_AXI_AWQOS_INT_M10
  `define AXI_AWQOS_INT_M10 `i_axi_AXI_AWQOS_INT_M10
`endif 

`ifdef i_axi_AXI_HAS_AWQOS_EXT_M11
  `define AXI_HAS_AWQOS_EXT_M11 `i_axi_AXI_HAS_AWQOS_EXT_M11
`endif 

`ifdef i_axi_AXI_AWQOS_EXT_M11
  `define AXI_AWQOS_EXT_M11 `i_axi_AXI_AWQOS_EXT_M11
`endif 

`ifdef i_axi_AXI_AWQOS_INT_M11
  `define AXI_AWQOS_INT_M11 `i_axi_AXI_AWQOS_INT_M11
`endif 

`ifdef i_axi_AXI_HAS_AWQOS_EXT_M12
  `define AXI_HAS_AWQOS_EXT_M12 `i_axi_AXI_HAS_AWQOS_EXT_M12
`endif 

`ifdef i_axi_AXI_AWQOS_EXT_M12
  `define AXI_AWQOS_EXT_M12 `i_axi_AXI_AWQOS_EXT_M12
`endif 

`ifdef i_axi_AXI_AWQOS_INT_M12
  `define AXI_AWQOS_INT_M12 `i_axi_AXI_AWQOS_INT_M12
`endif 

`ifdef i_axi_AXI_HAS_AWQOS_EXT_M13
  `define AXI_HAS_AWQOS_EXT_M13 `i_axi_AXI_HAS_AWQOS_EXT_M13
`endif 

`ifdef i_axi_AXI_AWQOS_EXT_M13
  `define AXI_AWQOS_EXT_M13 `i_axi_AXI_AWQOS_EXT_M13
`endif 

`ifdef i_axi_AXI_AWQOS_INT_M13
  `define AXI_AWQOS_INT_M13 `i_axi_AXI_AWQOS_INT_M13
`endif 

`ifdef i_axi_AXI_HAS_AWQOS_EXT_M14
  `define AXI_HAS_AWQOS_EXT_M14 `i_axi_AXI_HAS_AWQOS_EXT_M14
`endif 

`ifdef i_axi_AXI_AWQOS_EXT_M14
  `define AXI_AWQOS_EXT_M14 `i_axi_AXI_AWQOS_EXT_M14
`endif 

`ifdef i_axi_AXI_AWQOS_INT_M14
  `define AXI_AWQOS_INT_M14 `i_axi_AXI_AWQOS_INT_M14
`endif 

`ifdef i_axi_AXI_HAS_AWQOS_EXT_M15
  `define AXI_HAS_AWQOS_EXT_M15 `i_axi_AXI_HAS_AWQOS_EXT_M15
`endif 

`ifdef i_axi_AXI_AWQOS_EXT_M15
  `define AXI_AWQOS_EXT_M15 `i_axi_AXI_AWQOS_EXT_M15
`endif 

`ifdef i_axi_AXI_AWQOS_INT_M15
  `define AXI_AWQOS_INT_M15 `i_axi_AXI_AWQOS_INT_M15
`endif 

`ifdef i_axi_AXI_HAS_AWQOS_EXT_M16
  `define AXI_HAS_AWQOS_EXT_M16 `i_axi_AXI_HAS_AWQOS_EXT_M16
`endif 

`ifdef i_axi_AXI_AWQOS_EXT_M16
  `define AXI_AWQOS_EXT_M16 `i_axi_AXI_AWQOS_EXT_M16
`endif 

`ifdef i_axi_AXI_AWQOS_INT_M16
  `define AXI_AWQOS_INT_M16 `i_axi_AXI_AWQOS_INT_M16
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S0
  `define AXI_HAS_QOS_ARB_TYPE_ON_AR_S0 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S0
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S1
  `define AXI_HAS_QOS_ARB_TYPE_ON_AR_S1 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S1
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S2
  `define AXI_HAS_QOS_ARB_TYPE_ON_AR_S2 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S2
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S3
  `define AXI_HAS_QOS_ARB_TYPE_ON_AR_S3 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S3
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S4
  `define AXI_HAS_QOS_ARB_TYPE_ON_AR_S4 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S4
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S5
  `define AXI_HAS_QOS_ARB_TYPE_ON_AR_S5 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S5
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S6
  `define AXI_HAS_QOS_ARB_TYPE_ON_AR_S6 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S6
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S7
  `define AXI_HAS_QOS_ARB_TYPE_ON_AR_S7 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S7
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S8
  `define AXI_HAS_QOS_ARB_TYPE_ON_AR_S8 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S8
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S9
  `define AXI_HAS_QOS_ARB_TYPE_ON_AR_S9 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S9
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S10
  `define AXI_HAS_QOS_ARB_TYPE_ON_AR_S10 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S10
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S11
  `define AXI_HAS_QOS_ARB_TYPE_ON_AR_S11 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S11
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S12
  `define AXI_HAS_QOS_ARB_TYPE_ON_AR_S12 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S12
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S13
  `define AXI_HAS_QOS_ARB_TYPE_ON_AR_S13 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S13
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S14
  `define AXI_HAS_QOS_ARB_TYPE_ON_AR_S14 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S14
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S15
  `define AXI_HAS_QOS_ARB_TYPE_ON_AR_S15 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S15
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S16
  `define AXI_HAS_QOS_ARB_TYPE_ON_AR_S16 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AR_S16
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S0
  `define AXI_HAS_QOS_ARB_TYPE_ON_AW_S0 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S0
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S1
  `define AXI_HAS_QOS_ARB_TYPE_ON_AW_S1 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S1
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S2
  `define AXI_HAS_QOS_ARB_TYPE_ON_AW_S2 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S2
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S3
  `define AXI_HAS_QOS_ARB_TYPE_ON_AW_S3 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S3
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S4
  `define AXI_HAS_QOS_ARB_TYPE_ON_AW_S4 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S4
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S5
  `define AXI_HAS_QOS_ARB_TYPE_ON_AW_S5 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S5
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S6
  `define AXI_HAS_QOS_ARB_TYPE_ON_AW_S6 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S6
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S7
  `define AXI_HAS_QOS_ARB_TYPE_ON_AW_S7 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S7
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S8
  `define AXI_HAS_QOS_ARB_TYPE_ON_AW_S8 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S8
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S9
  `define AXI_HAS_QOS_ARB_TYPE_ON_AW_S9 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S9
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S10
  `define AXI_HAS_QOS_ARB_TYPE_ON_AW_S10 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S10
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S11
  `define AXI_HAS_QOS_ARB_TYPE_ON_AW_S11 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S11
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S12
  `define AXI_HAS_QOS_ARB_TYPE_ON_AW_S12 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S12
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S13
  `define AXI_HAS_QOS_ARB_TYPE_ON_AW_S13 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S13
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S14
  `define AXI_HAS_QOS_ARB_TYPE_ON_AW_S14 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S14
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S15
  `define AXI_HAS_QOS_ARB_TYPE_ON_AW_S15 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S15
`endif 

`ifdef i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S16
  `define AXI_HAS_QOS_ARB_TYPE_ON_AW_S16 `i_axi_AXI_HAS_QOS_ARB_TYPE_ON_AW_S16
`endif 

`ifdef i_axi_SNPS_RCE_INTERNAL_ON
  `define SNPS_RCE_INTERNAL_ON `i_axi_SNPS_RCE_INTERNAL_ON
`endif 

`ifdef i_axi_AXI_DW_GT_64
  `define AXI_DW_GT_64 `i_axi_AXI_DW_GT_64
`endif 

`ifdef i_axi_AXI_HAS_APB
  `define AXI_HAS_APB `i_axi_AXI_HAS_APB
`endif 

`ifdef i_axi_AXI_HAS_APB3
  `define AXI_HAS_APB3 `i_axi_AXI_HAS_APB3
`endif 

`ifdef i_axi_AXI_APB3
  `define AXI_APB3 `i_axi_AXI_APB3
`endif 

`ifdef i_axi_APB_DATA_WIDTH
  `define APB_DATA_WIDTH `i_axi_APB_DATA_WIDTH
`endif 

`ifdef i_axi_AXI_IC_REG_BASE_ADDR
  `define AXI_IC_REG_BASE_ADDR `i_axi_AXI_IC_REG_BASE_ADDR
`endif 

`ifdef i_axi_AXI_NUM_SYNC_FF
  `define AXI_NUM_SYNC_FF `i_axi_AXI_NUM_SYNC_FF
`endif 

`ifdef i_axi_DW_AXI_VERSION_ID
  `define DW_AXI_VERSION_ID `i_axi_DW_AXI_VERSION_ID
`endif 

`ifdef i_axi_AXI_VERIF_EN
  `define AXI_VERIF_EN `i_axi_AXI_VERIF_EN
`endif 

`ifdef i_axi_AXI_4
  `define AXI_4 `i_axi_AXI_4
`endif 

`ifdef i_axi_AXI_ACELITE
  `define AXI_ACELITE `i_axi_AXI_ACELITE
`endif 

`ifdef i_axi_AXI_HAS_REGIONS_S1
  `define AXI_HAS_REGIONS_S1 `i_axi_AXI_HAS_REGIONS_S1
`endif 

`ifdef i_axi_AXI_REGIONS_S1
  `define AXI_REGIONS_S1 `i_axi_AXI_REGIONS_S1
`endif 

`ifdef i_axi_AXI_HAS_REGIONS_S2
  `define AXI_HAS_REGIONS_S2 `i_axi_AXI_HAS_REGIONS_S2
`endif 

`ifdef i_axi_AXI_REGIONS_S2
  `define AXI_REGIONS_S2 `i_axi_AXI_REGIONS_S2
`endif 

`ifdef i_axi_AXI_HAS_REGIONS_S3
  `define AXI_HAS_REGIONS_S3 `i_axi_AXI_HAS_REGIONS_S3
`endif 

`ifdef i_axi_AXI_REGIONS_S3
  `define AXI_REGIONS_S3 `i_axi_AXI_REGIONS_S3
`endif 

`ifdef i_axi_AXI_HAS_REGIONS_S4
  `define AXI_HAS_REGIONS_S4 `i_axi_AXI_HAS_REGIONS_S4
`endif 

`ifdef i_axi_AXI_REGIONS_S4
  `define AXI_REGIONS_S4 `i_axi_AXI_REGIONS_S4
`endif 

`ifdef i_axi_AXI_HAS_REGIONS_S5
  `define AXI_HAS_REGIONS_S5 `i_axi_AXI_HAS_REGIONS_S5
`endif 

`ifdef i_axi_AXI_REGIONS_S5
  `define AXI_REGIONS_S5 `i_axi_AXI_REGIONS_S5
`endif 

`ifdef i_axi_AXI_HAS_REGIONS_S6
  `define AXI_HAS_REGIONS_S6 `i_axi_AXI_HAS_REGIONS_S6
`endif 

`ifdef i_axi_AXI_REGIONS_S6
  `define AXI_REGIONS_S6 `i_axi_AXI_REGIONS_S6
`endif 

`ifdef i_axi_AXI_HAS_REGIONS_S7
  `define AXI_HAS_REGIONS_S7 `i_axi_AXI_HAS_REGIONS_S7
`endif 

`ifdef i_axi_AXI_REGIONS_S7
  `define AXI_REGIONS_S7 `i_axi_AXI_REGIONS_S7
`endif 

`ifdef i_axi_AXI_HAS_REGIONS_S8
  `define AXI_HAS_REGIONS_S8 `i_axi_AXI_HAS_REGIONS_S8
`endif 

`ifdef i_axi_AXI_REGIONS_S8
  `define AXI_REGIONS_S8 `i_axi_AXI_REGIONS_S8
`endif 

`ifdef i_axi_AXI_HAS_REGIONS_S9
  `define AXI_HAS_REGIONS_S9 `i_axi_AXI_HAS_REGIONS_S9
`endif 

`ifdef i_axi_AXI_REGIONS_S9
  `define AXI_REGIONS_S9 `i_axi_AXI_REGIONS_S9
`endif 

`ifdef i_axi_AXI_HAS_REGIONS_S10
  `define AXI_HAS_REGIONS_S10 `i_axi_AXI_HAS_REGIONS_S10
`endif 

`ifdef i_axi_AXI_REGIONS_S10
  `define AXI_REGIONS_S10 `i_axi_AXI_REGIONS_S10
`endif 

`ifdef i_axi_AXI_HAS_REGIONS_S11
  `define AXI_HAS_REGIONS_S11 `i_axi_AXI_HAS_REGIONS_S11
`endif 

`ifdef i_axi_AXI_REGIONS_S11
  `define AXI_REGIONS_S11 `i_axi_AXI_REGIONS_S11
`endif 

`ifdef i_axi_AXI_HAS_REGIONS_S12
  `define AXI_HAS_REGIONS_S12 `i_axi_AXI_HAS_REGIONS_S12
`endif 

`ifdef i_axi_AXI_REGIONS_S12
  `define AXI_REGIONS_S12 `i_axi_AXI_REGIONS_S12
`endif 

`ifdef i_axi_AXI_HAS_REGIONS_S13
  `define AXI_HAS_REGIONS_S13 `i_axi_AXI_HAS_REGIONS_S13
`endif 

`ifdef i_axi_AXI_REGIONS_S13
  `define AXI_REGIONS_S13 `i_axi_AXI_REGIONS_S13
`endif 

`ifdef i_axi_AXI_HAS_REGIONS_S14
  `define AXI_HAS_REGIONS_S14 `i_axi_AXI_HAS_REGIONS_S14
`endif 

`ifdef i_axi_AXI_REGIONS_S14
  `define AXI_REGIONS_S14 `i_axi_AXI_REGIONS_S14
`endif 

`ifdef i_axi_AXI_HAS_REGIONS_S15
  `define AXI_HAS_REGIONS_S15 `i_axi_AXI_HAS_REGIONS_S15
`endif 

`ifdef i_axi_AXI_REGIONS_S15
  `define AXI_REGIONS_S15 `i_axi_AXI_REGIONS_S15
`endif 

`ifdef i_axi_AXI_HAS_REGIONS_S16
  `define AXI_HAS_REGIONS_S16 `i_axi_AXI_HAS_REGIONS_S16
`endif 

`ifdef i_axi_AXI_REGIONS_S16
  `define AXI_REGIONS_S16 `i_axi_AXI_REGIONS_S16
`endif 

`ifdef i_axi_AXI_HAS_REGIONS
  `define AXI_HAS_REGIONS `i_axi_AXI_HAS_REGIONS
`endif 

`ifdef i_axi_AXI_REGIONS
  `define AXI_REGIONS `i_axi_AXI_REGIONS
`endif 

`ifdef i_axi_AXI_LEGACY_LP_MODE
  `define AXI_LEGACY_LP_MODE `i_axi_AXI_LEGACY_LP_MODE
`endif 

`ifdef i_axi_AXI_BCM_TST_MODE
  `define AXI_BCM_TST_MODE `i_axi_AXI_BCM_TST_MODE
`endif 

`ifdef i_axi_AXI_BCM_CDC_INIT
  `define AXI_BCM_CDC_INIT `i_axi_AXI_BCM_CDC_INIT
`endif 

`ifdef i_axi_DWC_NO_TST_MODE
  `define DWC_NO_TST_MODE `i_axi_DWC_NO_TST_MODE
`endif 

`ifdef i_axi_DWC_NO_CDC_INIT
  `define DWC_NO_CDC_INIT `i_axi_DWC_NO_CDC_INIT
`endif 

`ifdef i_axi___GUARD__DW_AXI_CONSTANTS__VH__
  `define __GUARD__DW_AXI_CONSTANTS__VH__ `i_axi___GUARD__DW_AXI_CONSTANTS__VH__
`endif 

`ifdef i_axi_AXI_BSW
  `define AXI_BSW `i_axi_AXI_BSW
`endif 

`ifdef i_axi_AXI_BTW
  `define AXI_BTW `i_axi_AXI_BTW
`endif 

`ifdef i_axi_AXI_LTW
  `define AXI_LTW `i_axi_AXI_LTW
`endif 

`ifdef i_axi_AXI_CTW
  `define AXI_CTW `i_axi_AXI_CTW
`endif 

`ifdef i_axi_AXI_PTW
  `define AXI_PTW `i_axi_AXI_PTW
`endif 

`ifdef i_axi_AXI_BRW
  `define AXI_BRW `i_axi_AXI_BRW
`endif 

`ifdef i_axi_AXI_RRW
  `define AXI_RRW `i_axi_AXI_RRW
`endif 

`ifdef i_axi_AXI_SW
  `define AXI_SW `i_axi_AXI_SW
`endif 

`ifdef i_axi_AXI_MAX_NUM_MST_SLVS
  `define AXI_MAX_NUM_MST_SLVS `i_axi_AXI_MAX_NUM_MST_SLVS
`endif 

`ifdef i_axi_AXI_MAX_NUM_USR_MSTS
  `define AXI_MAX_NUM_USR_MSTS `i_axi_AXI_MAX_NUM_USR_MSTS
`endif 

`ifdef i_axi_AXI_MAX_NUM_USR_SLVS
  `define AXI_MAX_NUM_USR_SLVS `i_axi_AXI_MAX_NUM_USR_SLVS
`endif 

`ifdef i_axi_AXI_LT_NORM
  `define AXI_LT_NORM `i_axi_AXI_LT_NORM
`endif 

`ifdef i_axi_AXI_LT_EX
  `define AXI_LT_EX `i_axi_AXI_LT_EX
`endif 

`ifdef i_axi_AXI_LT_LOCK
  `define AXI_LT_LOCK `i_axi_AXI_LT_LOCK
`endif 

`ifdef i_axi_AXI_PT_PRVLGD
  `define AXI_PT_PRVLGD `i_axi_AXI_PT_PRVLGD
`endif 

`ifdef i_axi_AXI_PT_NORM
  `define AXI_PT_NORM `i_axi_AXI_PT_NORM
`endif 

`ifdef i_axi_AXI_PT_SECURE
  `define AXI_PT_SECURE `i_axi_AXI_PT_SECURE
`endif 

`ifdef i_axi_AXI_PT_NSECURE
  `define AXI_PT_NSECURE `i_axi_AXI_PT_NSECURE
`endif 

`ifdef i_axi_AXI_PT_INSTRUCT
  `define AXI_PT_INSTRUCT `i_axi_AXI_PT_INSTRUCT
`endif 

`ifdef i_axi_AXI_PT_DATA
  `define AXI_PT_DATA `i_axi_AXI_PT_DATA
`endif 

`ifdef i_axi_AXI_PT_PRVLGD_BIT
  `define AXI_PT_PRVLGD_BIT `i_axi_AXI_PT_PRVLGD_BIT
`endif 

`ifdef i_axi_AXI_PT_INSTRUCT_BIT
  `define AXI_PT_INSTRUCT_BIT `i_axi_AXI_PT_INSTRUCT_BIT
`endif 

`ifdef i_axi_AXI_RESP_OKAY
  `define AXI_RESP_OKAY `i_axi_AXI_RESP_OKAY
`endif 

`ifdef i_axi_AXI_RESP_EXOKAY
  `define AXI_RESP_EXOKAY `i_axi_AXI_RESP_EXOKAY
`endif 

`ifdef i_axi_AXI_RESP_SLVERR
  `define AXI_RESP_SLVERR `i_axi_AXI_RESP_SLVERR
`endif 

`ifdef i_axi_AXI_RESP_DECERR
  `define AXI_RESP_DECERR `i_axi_AXI_RESP_DECERR
`endif 

`ifdef i_axi_AXI_TMO_COMB
  `define AXI_TMO_COMB `i_axi_AXI_TMO_COMB
`endif 

`ifdef i_axi_AXI_TMO_FRWD
  `define AXI_TMO_FRWD `i_axi_AXI_TMO_FRWD
`endif 

`ifdef i_axi_AXI_TMO_FULL
  `define AXI_TMO_FULL `i_axi_AXI_TMO_FULL
`endif 

`ifdef i_axi_AXI_NOREQ_LOCKING
  `define AXI_NOREQ_LOCKING `i_axi_AXI_NOREQ_LOCKING
`endif 

`ifdef i_axi_AXI_REQ_LOCKING
  `define AXI_REQ_LOCKING `i_axi_AXI_REQ_LOCKING
`endif 

`ifdef i_axi_AXI_ARB_TYPE_DP
  `define AXI_ARB_TYPE_DP `i_axi_AXI_ARB_TYPE_DP
`endif 

`ifdef i_axi_AXI_ARB_TYPE_FCFS
  `define AXI_ARB_TYPE_FCFS `i_axi_AXI_ARB_TYPE_FCFS
`endif 

`ifdef i_axi_AXI_ARB_TYPE_2T
  `define AXI_ARB_TYPE_2T `i_axi_AXI_ARB_TYPE_2T
`endif 

`ifdef i_axi_AXI_ARB_TYPE_USER
  `define AXI_ARB_TYPE_USER `i_axi_AXI_ARB_TYPE_USER
`endif 

`ifdef i_axi_AXI_ARB_TYPE_QOS
  `define AXI_ARB_TYPE_QOS `i_axi_AXI_ARB_TYPE_QOS
`endif 

`ifdef i_axi_AXI_W_CH
  `define AXI_W_CH `i_axi_AXI_W_CH
`endif 

`ifdef i_axi_AXI_NOT_W_CH
  `define AXI_NOT_W_CH `i_axi_AXI_NOT_W_CH
`endif 

`ifdef i_axi_AXI_AW_CH
  `define AXI_AW_CH `i_axi_AXI_AW_CH
`endif 

`ifdef i_axi_AXI_NOT_AW_CH
  `define AXI_NOT_AW_CH `i_axi_AXI_NOT_AW_CH
`endif 

`ifdef i_axi_AXI_R_CH
  `define AXI_R_CH `i_axi_AXI_R_CH
`endif 

`ifdef i_axi_AXI_NOT_R_CH
  `define AXI_NOT_R_CH `i_axi_AXI_NOT_R_CH
`endif 

`ifdef i_axi_AXI_ADDR_CH
  `define AXI_ADDR_CH `i_axi_AXI_ADDR_CH
`endif 

`ifdef i_axi_AXI_NOT_ADDR_CH
  `define AXI_NOT_ADDR_CH `i_axi_AXI_NOT_ADDR_CH
`endif 

`ifdef i_axi_USE_INT_GI
  `define USE_INT_GI `i_axi_USE_INT_GI
`endif 

`ifdef i_axi_USE_EXT_GI
  `define USE_EXT_GI `i_axi_USE_EXT_GI
`endif 

`ifdef i_axi_AXI_SHARED
  `define AXI_SHARED `i_axi_AXI_SHARED
`endif 

`ifdef i_axi_AXI_NOT_SHARED
  `define AXI_NOT_SHARED `i_axi_AXI_NOT_SHARED
`endif 

`ifdef i_axi_AXI_HOLD_VLD_OTHER_S_W
  `define AXI_HOLD_VLD_OTHER_S_W `i_axi_AXI_HOLD_VLD_OTHER_S_W
`endif 

`ifdef i_axi_AXI_HOLD_VLD_OTHER_M_W
  `define AXI_HOLD_VLD_OTHER_M_W `i_axi_AXI_HOLD_VLD_OTHER_M_W
`endif 

`ifdef i_axi_AXI_ARPYLD_PROT_RHS
  `define AXI_ARPYLD_PROT_RHS `i_axi_AXI_ARPYLD_PROT_RHS
`endif 

`ifdef i_axi_AXI_ARPYLD_PROT_LHS
  `define AXI_ARPYLD_PROT_LHS `i_axi_AXI_ARPYLD_PROT_LHS
`endif 

`ifdef i_axi_AXI_ARPYLD_PROT
  `define AXI_ARPYLD_PROT `i_axi_AXI_ARPYLD_PROT
`endif 

`ifdef i_axi_AXI_ARPYLD_CACHE_RHS
  `define AXI_ARPYLD_CACHE_RHS `i_axi_AXI_ARPYLD_CACHE_RHS
`endif 

`ifdef i_axi_AXI_ARPYLD_CACHE_LHS
  `define AXI_ARPYLD_CACHE_LHS `i_axi_AXI_ARPYLD_CACHE_LHS
`endif 

`ifdef i_axi_AXI_ARPYLD_CACHE
  `define AXI_ARPYLD_CACHE `i_axi_AXI_ARPYLD_CACHE
`endif 

`ifdef i_axi_AXI_ARPYLD_LOCK_RHS
  `define AXI_ARPYLD_LOCK_RHS `i_axi_AXI_ARPYLD_LOCK_RHS
`endif 

`ifdef i_axi_AXI_ARPYLD_LOCK_LHS
  `define AXI_ARPYLD_LOCK_LHS `i_axi_AXI_ARPYLD_LOCK_LHS
`endif 

`ifdef i_axi_AXI_ARPYLD_LOCK
  `define AXI_ARPYLD_LOCK `i_axi_AXI_ARPYLD_LOCK
`endif 

`ifdef i_axi_AXI_ARPYLD_BURST_RHS
  `define AXI_ARPYLD_BURST_RHS `i_axi_AXI_ARPYLD_BURST_RHS
`endif 

`ifdef i_axi_AXI_ARPYLD_BURST_LHS
  `define AXI_ARPYLD_BURST_LHS `i_axi_AXI_ARPYLD_BURST_LHS
`endif 

`ifdef i_axi_AXI_ARPYLD_BURST
  `define AXI_ARPYLD_BURST `i_axi_AXI_ARPYLD_BURST
`endif 

`ifdef i_axi_AXI_ARPYLD_SIZE_RHS
  `define AXI_ARPYLD_SIZE_RHS `i_axi_AXI_ARPYLD_SIZE_RHS
`endif 

`ifdef i_axi_AXI_ARPYLD_SIZE_LHS
  `define AXI_ARPYLD_SIZE_LHS `i_axi_AXI_ARPYLD_SIZE_LHS
`endif 

`ifdef i_axi_AXI_ARPYLD_SIZE
  `define AXI_ARPYLD_SIZE `i_axi_AXI_ARPYLD_SIZE
`endif 

`ifdef i_axi_AXI_ARPYLD_LEN_RHS
  `define AXI_ARPYLD_LEN_RHS `i_axi_AXI_ARPYLD_LEN_RHS
`endif 

`ifdef i_axi_AXI_ARPYLD_LEN_LHS
  `define AXI_ARPYLD_LEN_LHS `i_axi_AXI_ARPYLD_LEN_LHS
`endif 

`ifdef i_axi_AXI_ARPYLD_LEN
  `define AXI_ARPYLD_LEN `i_axi_AXI_ARPYLD_LEN
`endif 

`ifdef i_axi_AXI_ARPYLD_ADDR_RHS
  `define AXI_ARPYLD_ADDR_RHS `i_axi_AXI_ARPYLD_ADDR_RHS
`endif 

`ifdef i_axi_AXI_ARPYLD_ADDR_LHS
  `define AXI_ARPYLD_ADDR_LHS `i_axi_AXI_ARPYLD_ADDR_LHS
`endif 

`ifdef i_axi_AXI_ARPYLD_ADDR
  `define AXI_ARPYLD_ADDR `i_axi_AXI_ARPYLD_ADDR
`endif 

`ifdef i_axi_AXI_ARPYLD_ID_RHS_M
  `define AXI_ARPYLD_ID_RHS_M `i_axi_AXI_ARPYLD_ID_RHS_M
`endif 

`ifdef i_axi_AXI_ARPYLD_ID_LHS_M
  `define AXI_ARPYLD_ID_LHS_M `i_axi_AXI_ARPYLD_ID_LHS_M
`endif 

`ifdef i_axi_AXI_ARPYLD_ID_M
  `define AXI_ARPYLD_ID_M `i_axi_AXI_ARPYLD_ID_M
`endif 

`ifdef i_axi_AXI_ARPYLD_ID_RHS_S
  `define AXI_ARPYLD_ID_RHS_S `i_axi_AXI_ARPYLD_ID_RHS_S
`endif 

`ifdef i_axi_AXI_ARPYLD_ID_LHS_S
  `define AXI_ARPYLD_ID_LHS_S `i_axi_AXI_ARPYLD_ID_LHS_S
`endif 

`ifdef i_axi_AXI_ARPYLD_ID_S
  `define AXI_ARPYLD_ID_S `i_axi_AXI_ARPYLD_ID_S
`endif 

`ifdef i_axi_AXI_RPYLD_LAST_LHS
  `define AXI_RPYLD_LAST_LHS `i_axi_AXI_RPYLD_LAST_LHS
`endif 

`ifdef i_axi_AXI_RPYLD_LAST
  `define AXI_RPYLD_LAST `i_axi_AXI_RPYLD_LAST
`endif 

`ifdef i_axi_AXI_RPYLD_RESP_RHS
  `define AXI_RPYLD_RESP_RHS `i_axi_AXI_RPYLD_RESP_RHS
`endif 

`ifdef i_axi_AXI_RPYLD_RESP_LHS
  `define AXI_RPYLD_RESP_LHS `i_axi_AXI_RPYLD_RESP_LHS
`endif 

`ifdef i_axi_AXI_RPYLD_RESP
  `define AXI_RPYLD_RESP `i_axi_AXI_RPYLD_RESP
`endif 

`ifdef i_axi_AXI_RPYLD_DATA_RHS
  `define AXI_RPYLD_DATA_RHS `i_axi_AXI_RPYLD_DATA_RHS
`endif 

`ifdef i_axi_AXI_RPYLD_DATA_LHS
  `define AXI_RPYLD_DATA_LHS `i_axi_AXI_RPYLD_DATA_LHS
`endif 

`ifdef i_axi_AXI_RPYLD_DATA
  `define AXI_RPYLD_DATA `i_axi_AXI_RPYLD_DATA
`endif 

`ifdef i_axi_AXI_RPYLD_ID_RHS_M
  `define AXI_RPYLD_ID_RHS_M `i_axi_AXI_RPYLD_ID_RHS_M
`endif 

`ifdef i_axi_AXI_RPYLD_ID_LHS_M
  `define AXI_RPYLD_ID_LHS_M `i_axi_AXI_RPYLD_ID_LHS_M
`endif 

`ifdef i_axi_AXI_RPYLD_ID_M
  `define AXI_RPYLD_ID_M `i_axi_AXI_RPYLD_ID_M
`endif 

`ifdef i_axi_AXI_RPYLD_ID_RHS_S
  `define AXI_RPYLD_ID_RHS_S `i_axi_AXI_RPYLD_ID_RHS_S
`endif 

`ifdef i_axi_AXI_RPYLD_ID_LHS_S
  `define AXI_RPYLD_ID_LHS_S `i_axi_AXI_RPYLD_ID_LHS_S
`endif 

`ifdef i_axi_AXI_RPYLD_ID_S
  `define AXI_RPYLD_ID_S `i_axi_AXI_RPYLD_ID_S
`endif 

`ifdef i_axi_AXI_AWPYLD_PROT_RHS
  `define AXI_AWPYLD_PROT_RHS `i_axi_AXI_AWPYLD_PROT_RHS
`endif 

`ifdef i_axi_AXI_AWPYLD_PROT_LHS
  `define AXI_AWPYLD_PROT_LHS `i_axi_AXI_AWPYLD_PROT_LHS
`endif 

`ifdef i_axi_AXI_AWPYLD_PROT
  `define AXI_AWPYLD_PROT `i_axi_AXI_AWPYLD_PROT
`endif 

`ifdef i_axi_AXI_AWPYLD_CACHE_RHS
  `define AXI_AWPYLD_CACHE_RHS `i_axi_AXI_AWPYLD_CACHE_RHS
`endif 

`ifdef i_axi_AXI_AWPYLD_CACHE_LHS
  `define AXI_AWPYLD_CACHE_LHS `i_axi_AXI_AWPYLD_CACHE_LHS
`endif 

`ifdef i_axi_AXI_AWPYLD_CACHE
  `define AXI_AWPYLD_CACHE `i_axi_AXI_AWPYLD_CACHE
`endif 

`ifdef i_axi_AXI_AWPYLD_LOCK_RHS
  `define AXI_AWPYLD_LOCK_RHS `i_axi_AXI_AWPYLD_LOCK_RHS
`endif 

`ifdef i_axi_AXI_AWPYLD_LOCK_LHS
  `define AXI_AWPYLD_LOCK_LHS `i_axi_AXI_AWPYLD_LOCK_LHS
`endif 

`ifdef i_axi_AXI_AWPYLD_LOCK
  `define AXI_AWPYLD_LOCK `i_axi_AXI_AWPYLD_LOCK
`endif 

`ifdef i_axi_AXI_AWPYLD_BURST_RHS
  `define AXI_AWPYLD_BURST_RHS `i_axi_AXI_AWPYLD_BURST_RHS
`endif 

`ifdef i_axi_AXI_AWPYLD_BURST_LHS
  `define AXI_AWPYLD_BURST_LHS `i_axi_AXI_AWPYLD_BURST_LHS
`endif 

`ifdef i_axi_AXI_AWPYLD_BURST
  `define AXI_AWPYLD_BURST `i_axi_AXI_AWPYLD_BURST
`endif 

`ifdef i_axi_AXI_AWPYLD_SIZE_RHS
  `define AXI_AWPYLD_SIZE_RHS `i_axi_AXI_AWPYLD_SIZE_RHS
`endif 

`ifdef i_axi_AXI_AWPYLD_SIZE_LHS
  `define AXI_AWPYLD_SIZE_LHS `i_axi_AXI_AWPYLD_SIZE_LHS
`endif 

`ifdef i_axi_AXI_AWPYLD_SIZE
  `define AXI_AWPYLD_SIZE `i_axi_AXI_AWPYLD_SIZE
`endif 

`ifdef i_axi_AXI_AWPYLD_LEN_RHS
  `define AXI_AWPYLD_LEN_RHS `i_axi_AXI_AWPYLD_LEN_RHS
`endif 

`ifdef i_axi_AXI_AWPYLD_LEN_LHS
  `define AXI_AWPYLD_LEN_LHS `i_axi_AXI_AWPYLD_LEN_LHS
`endif 

`ifdef i_axi_AXI_AWPYLD_LEN
  `define AXI_AWPYLD_LEN `i_axi_AXI_AWPYLD_LEN
`endif 

`ifdef i_axi_AXI_AWPYLD_ADDR_RHS
  `define AXI_AWPYLD_ADDR_RHS `i_axi_AXI_AWPYLD_ADDR_RHS
`endif 

`ifdef i_axi_AXI_AWPYLD_ADDR_LHS
  `define AXI_AWPYLD_ADDR_LHS `i_axi_AXI_AWPYLD_ADDR_LHS
`endif 

`ifdef i_axi_AXI_AWPYLD_ADDR
  `define AXI_AWPYLD_ADDR `i_axi_AXI_AWPYLD_ADDR
`endif 

`ifdef i_axi_AXI_AWPYLD_ID_RHS_M
  `define AXI_AWPYLD_ID_RHS_M `i_axi_AXI_AWPYLD_ID_RHS_M
`endif 

`ifdef i_axi_AXI_AWPYLD_ID_LHS_M
  `define AXI_AWPYLD_ID_LHS_M `i_axi_AXI_AWPYLD_ID_LHS_M
`endif 

`ifdef i_axi_AXI_AWPYLD_ID_M
  `define AXI_AWPYLD_ID_M `i_axi_AXI_AWPYLD_ID_M
`endif 

`ifdef i_axi_AXI_AWPYLD_ID_RHS_S
  `define AXI_AWPYLD_ID_RHS_S `i_axi_AXI_AWPYLD_ID_RHS_S
`endif 

`ifdef i_axi_AXI_AWPYLD_ID_LHS_S
  `define AXI_AWPYLD_ID_LHS_S `i_axi_AXI_AWPYLD_ID_LHS_S
`endif 

`ifdef i_axi_AXI_AWPYLD_ID_S
  `define AXI_AWPYLD_ID_S `i_axi_AXI_AWPYLD_ID_S
`endif 

`ifdef i_axi_AXI_WPYLD_LAST_LHS
  `define AXI_WPYLD_LAST_LHS `i_axi_AXI_WPYLD_LAST_LHS
`endif 

`ifdef i_axi_AXI_WPYLD_LAST
  `define AXI_WPYLD_LAST `i_axi_AXI_WPYLD_LAST
`endif 

`ifdef i_axi_AXI_WPYLD_STRB_RHS
  `define AXI_WPYLD_STRB_RHS `i_axi_AXI_WPYLD_STRB_RHS
`endif 

`ifdef i_axi_AXI_WPYLD_STRB_LHS
  `define AXI_WPYLD_STRB_LHS `i_axi_AXI_WPYLD_STRB_LHS
`endif 

`ifdef i_axi_AXI_WPYLD_STRB
  `define AXI_WPYLD_STRB `i_axi_AXI_WPYLD_STRB
`endif 

`ifdef i_axi_AXI_WPYLD_DATA_RHS
  `define AXI_WPYLD_DATA_RHS `i_axi_AXI_WPYLD_DATA_RHS
`endif 

`ifdef i_axi_AXI_WPYLD_DATA_LHS
  `define AXI_WPYLD_DATA_LHS `i_axi_AXI_WPYLD_DATA_LHS
`endif 

`ifdef i_axi_AXI_WPYLD_DATA
  `define AXI_WPYLD_DATA `i_axi_AXI_WPYLD_DATA
`endif 

`ifdef i_axi_AXI_WPYLD_ID_RHS_M
  `define AXI_WPYLD_ID_RHS_M `i_axi_AXI_WPYLD_ID_RHS_M
`endif 

`ifdef i_axi_AXI_WPYLD_ID_LHS_M
  `define AXI_WPYLD_ID_LHS_M `i_axi_AXI_WPYLD_ID_LHS_M
`endif 

`ifdef i_axi_AXI_WPYLD_ID_M
  `define AXI_WPYLD_ID_M `i_axi_AXI_WPYLD_ID_M
`endif 

`ifdef i_axi_AXI_WPYLD_ID_RHS_S
  `define AXI_WPYLD_ID_RHS_S `i_axi_AXI_WPYLD_ID_RHS_S
`endif 

`ifdef i_axi_AXI_WPYLD_ID_LHS_S
  `define AXI_WPYLD_ID_LHS_S `i_axi_AXI_WPYLD_ID_LHS_S
`endif 

`ifdef i_axi_AXI_WPYLD_ID_S
  `define AXI_WPYLD_ID_S `i_axi_AXI_WPYLD_ID_S
`endif 

`ifdef i_axi_AXI_BPYLD_RESP_RHS
  `define AXI_BPYLD_RESP_RHS `i_axi_AXI_BPYLD_RESP_RHS
`endif 

`ifdef i_axi_AXI_BPYLD_RESP_LHS
  `define AXI_BPYLD_RESP_LHS `i_axi_AXI_BPYLD_RESP_LHS
`endif 

`ifdef i_axi_AXI_BPYLD_RESP
  `define AXI_BPYLD_RESP `i_axi_AXI_BPYLD_RESP
`endif 

`ifdef i_axi_AXI_BPYLD_ID_RHS_M
  `define AXI_BPYLD_ID_RHS_M `i_axi_AXI_BPYLD_ID_RHS_M
`endif 

`ifdef i_axi_AXI_BPYLD_ID_LHS_M
  `define AXI_BPYLD_ID_LHS_M `i_axi_AXI_BPYLD_ID_LHS_M
`endif 

`ifdef i_axi_AXI_BPYLD_ID_M
  `define AXI_BPYLD_ID_M `i_axi_AXI_BPYLD_ID_M
`endif 

`ifdef i_axi_AXI_BPYLD_ID_RHS_S
  `define AXI_BPYLD_ID_RHS_S `i_axi_AXI_BPYLD_ID_RHS_S
`endif 

`ifdef i_axi_AXI_BPYLD_ID_LHS_S
  `define AXI_BPYLD_ID_LHS_S `i_axi_AXI_BPYLD_ID_LHS_S
`endif 

`ifdef i_axi_AXI_BPYLD_ID_S
  `define AXI_BPYLD_ID_S `i_axi_AXI_BPYLD_ID_S
`endif 

`ifdef i_axi_AXI_QOSW
  `define AXI_QOSW `i_axi_AXI_QOSW
`endif 

`ifdef i_axi_IC_ADDR_SLICE_LHS
  `define IC_ADDR_SLICE_LHS `i_axi_IC_ADDR_SLICE_LHS
`endif 

`ifdef i_axi_MAX_APB_DATA_WIDTH
  `define MAX_APB_DATA_WIDTH `i_axi_MAX_APB_DATA_WIDTH
`endif 

`ifdef i_axi_REG_XCT_RATE_W
  `define REG_XCT_RATE_W `i_axi_REG_XCT_RATE_W
`endif 

`ifdef i_axi_REG_BURSTINESS_W
  `define REG_BURSTINESS_W `i_axi_REG_BURSTINESS_W
`endif 

`ifdef i_axi_REG_PEAK_RATE_W
  `define REG_PEAK_RATE_W `i_axi_REG_PEAK_RATE_W
`endif 

`ifdef i_axi_APB_ADDR_WIDTH
  `define APB_ADDR_WIDTH `i_axi_APB_ADDR_WIDTH
`endif 

`ifdef i_axi_AXI_ALSW
  `define AXI_ALSW `i_axi_AXI_ALSW
`endif 

`ifdef i_axi_AXI_ALDW
  `define AXI_ALDW `i_axi_AXI_ALDW
`endif 

`ifdef i_axi_AXI_ALBW
  `define AXI_ALBW `i_axi_AXI_ALBW
`endif 

`ifdef i_axi_AXI_REGIONW
  `define AXI_REGIONW `i_axi_AXI_REGIONW
`endif 

`ifdef i_axi_PL_BUF_AW
  `define PL_BUF_AW `i_axi_PL_BUF_AW
`endif 

`ifdef i_axi_PL_BUF_AR
  `define PL_BUF_AR `i_axi_PL_BUF_AR
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AW_M1
  `define ACT_ID_BUF_POINTER_W_AW_M1 `i_axi_ACT_ID_BUF_POINTER_W_AW_M1
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M1
  `define LOG2_ACT_ID_BUF_POINTER_W_AW_M1 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M1
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AR_M1
  `define ACT_ID_BUF_POINTER_W_AR_M1 `i_axi_ACT_ID_BUF_POINTER_W_AR_M1
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M1
  `define LOG2_ACT_ID_BUF_POINTER_W_AR_M1 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M1
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AW_M2
  `define ACT_ID_BUF_POINTER_W_AW_M2 `i_axi_ACT_ID_BUF_POINTER_W_AW_M2
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M2
  `define LOG2_ACT_ID_BUF_POINTER_W_AW_M2 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M2
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AR_M2
  `define ACT_ID_BUF_POINTER_W_AR_M2 `i_axi_ACT_ID_BUF_POINTER_W_AR_M2
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M2
  `define LOG2_ACT_ID_BUF_POINTER_W_AR_M2 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M2
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AW_M3
  `define ACT_ID_BUF_POINTER_W_AW_M3 `i_axi_ACT_ID_BUF_POINTER_W_AW_M3
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M3
  `define LOG2_ACT_ID_BUF_POINTER_W_AW_M3 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M3
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AR_M3
  `define ACT_ID_BUF_POINTER_W_AR_M3 `i_axi_ACT_ID_BUF_POINTER_W_AR_M3
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M3
  `define LOG2_ACT_ID_BUF_POINTER_W_AR_M3 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M3
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AW_M4
  `define ACT_ID_BUF_POINTER_W_AW_M4 `i_axi_ACT_ID_BUF_POINTER_W_AW_M4
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M4
  `define LOG2_ACT_ID_BUF_POINTER_W_AW_M4 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M4
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AR_M4
  `define ACT_ID_BUF_POINTER_W_AR_M4 `i_axi_ACT_ID_BUF_POINTER_W_AR_M4
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M4
  `define LOG2_ACT_ID_BUF_POINTER_W_AR_M4 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M4
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AW_M5
  `define ACT_ID_BUF_POINTER_W_AW_M5 `i_axi_ACT_ID_BUF_POINTER_W_AW_M5
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M5
  `define LOG2_ACT_ID_BUF_POINTER_W_AW_M5 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M5
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AR_M5
  `define ACT_ID_BUF_POINTER_W_AR_M5 `i_axi_ACT_ID_BUF_POINTER_W_AR_M5
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M5
  `define LOG2_ACT_ID_BUF_POINTER_W_AR_M5 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M5
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AW_M6
  `define ACT_ID_BUF_POINTER_W_AW_M6 `i_axi_ACT_ID_BUF_POINTER_W_AW_M6
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M6
  `define LOG2_ACT_ID_BUF_POINTER_W_AW_M6 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M6
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AR_M6
  `define ACT_ID_BUF_POINTER_W_AR_M6 `i_axi_ACT_ID_BUF_POINTER_W_AR_M6
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M6
  `define LOG2_ACT_ID_BUF_POINTER_W_AR_M6 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M6
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AW_M7
  `define ACT_ID_BUF_POINTER_W_AW_M7 `i_axi_ACT_ID_BUF_POINTER_W_AW_M7
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M7
  `define LOG2_ACT_ID_BUF_POINTER_W_AW_M7 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M7
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AR_M7
  `define ACT_ID_BUF_POINTER_W_AR_M7 `i_axi_ACT_ID_BUF_POINTER_W_AR_M7
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M7
  `define LOG2_ACT_ID_BUF_POINTER_W_AR_M7 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M7
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AW_M8
  `define ACT_ID_BUF_POINTER_W_AW_M8 `i_axi_ACT_ID_BUF_POINTER_W_AW_M8
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M8
  `define LOG2_ACT_ID_BUF_POINTER_W_AW_M8 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M8
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AR_M8
  `define ACT_ID_BUF_POINTER_W_AR_M8 `i_axi_ACT_ID_BUF_POINTER_W_AR_M8
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M8
  `define LOG2_ACT_ID_BUF_POINTER_W_AR_M8 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M8
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AW_M9
  `define ACT_ID_BUF_POINTER_W_AW_M9 `i_axi_ACT_ID_BUF_POINTER_W_AW_M9
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M9
  `define LOG2_ACT_ID_BUF_POINTER_W_AW_M9 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M9
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AR_M9
  `define ACT_ID_BUF_POINTER_W_AR_M9 `i_axi_ACT_ID_BUF_POINTER_W_AR_M9
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M9
  `define LOG2_ACT_ID_BUF_POINTER_W_AR_M9 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M9
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AW_M10
  `define ACT_ID_BUF_POINTER_W_AW_M10 `i_axi_ACT_ID_BUF_POINTER_W_AW_M10
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M10
  `define LOG2_ACT_ID_BUF_POINTER_W_AW_M10 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M10
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AR_M10
  `define ACT_ID_BUF_POINTER_W_AR_M10 `i_axi_ACT_ID_BUF_POINTER_W_AR_M10
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M10
  `define LOG2_ACT_ID_BUF_POINTER_W_AR_M10 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M10
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AW_M11
  `define ACT_ID_BUF_POINTER_W_AW_M11 `i_axi_ACT_ID_BUF_POINTER_W_AW_M11
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M11
  `define LOG2_ACT_ID_BUF_POINTER_W_AW_M11 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M11
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AR_M11
  `define ACT_ID_BUF_POINTER_W_AR_M11 `i_axi_ACT_ID_BUF_POINTER_W_AR_M11
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M11
  `define LOG2_ACT_ID_BUF_POINTER_W_AR_M11 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M11
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AW_M12
  `define ACT_ID_BUF_POINTER_W_AW_M12 `i_axi_ACT_ID_BUF_POINTER_W_AW_M12
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M12
  `define LOG2_ACT_ID_BUF_POINTER_W_AW_M12 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M12
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AR_M12
  `define ACT_ID_BUF_POINTER_W_AR_M12 `i_axi_ACT_ID_BUF_POINTER_W_AR_M12
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M12
  `define LOG2_ACT_ID_BUF_POINTER_W_AR_M12 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M12
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AW_M13
  `define ACT_ID_BUF_POINTER_W_AW_M13 `i_axi_ACT_ID_BUF_POINTER_W_AW_M13
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M13
  `define LOG2_ACT_ID_BUF_POINTER_W_AW_M13 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M13
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AR_M13
  `define ACT_ID_BUF_POINTER_W_AR_M13 `i_axi_ACT_ID_BUF_POINTER_W_AR_M13
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M13
  `define LOG2_ACT_ID_BUF_POINTER_W_AR_M13 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M13
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AW_M14
  `define ACT_ID_BUF_POINTER_W_AW_M14 `i_axi_ACT_ID_BUF_POINTER_W_AW_M14
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M14
  `define LOG2_ACT_ID_BUF_POINTER_W_AW_M14 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M14
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AR_M14
  `define ACT_ID_BUF_POINTER_W_AR_M14 `i_axi_ACT_ID_BUF_POINTER_W_AR_M14
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M14
  `define LOG2_ACT_ID_BUF_POINTER_W_AR_M14 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M14
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AW_M15
  `define ACT_ID_BUF_POINTER_W_AW_M15 `i_axi_ACT_ID_BUF_POINTER_W_AW_M15
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M15
  `define LOG2_ACT_ID_BUF_POINTER_W_AW_M15 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M15
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AR_M15
  `define ACT_ID_BUF_POINTER_W_AR_M15 `i_axi_ACT_ID_BUF_POINTER_W_AR_M15
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M15
  `define LOG2_ACT_ID_BUF_POINTER_W_AR_M15 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M15
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AW_M16
  `define ACT_ID_BUF_POINTER_W_AW_M16 `i_axi_ACT_ID_BUF_POINTER_W_AW_M16
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M16
  `define LOG2_ACT_ID_BUF_POINTER_W_AW_M16 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AW_M16
`endif 

`ifdef i_axi_ACT_ID_BUF_POINTER_W_AR_M16
  `define ACT_ID_BUF_POINTER_W_AR_M16 `i_axi_ACT_ID_BUF_POINTER_W_AR_M16
`endif 

`ifdef i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M16
  `define LOG2_ACT_ID_BUF_POINTER_W_AR_M16 `i_axi_LOG2_ACT_ID_BUF_POINTER_W_AR_M16
`endif 

`ifdef i_axi_AXI_HAS_WID
  `define AXI_HAS_WID `i_axi_AXI_HAS_WID
`endif 

`ifdef i_axi___GUARD__DW_AXI_BCM_PARAMS__VH__
  `define __GUARD__DW_AXI_BCM_PARAMS__VH__ `i_axi___GUARD__DW_AXI_BCM_PARAMS__VH__
`endif 

`ifdef i_axi_DW_AXI_RM_BCM00_AND
  `define DW_AXI_RM_BCM00_AND `i_axi_DW_AXI_RM_BCM00_AND
`endif 

`ifdef i_axi_DW_AXI_RM_BCM00_ATPG_MX
  `define DW_AXI_RM_BCM00_ATPG_MX `i_axi_DW_AXI_RM_BCM00_ATPG_MX
`endif 

`ifdef i_axi_DW_AXI_RM_BCM00_CK_AND
  `define DW_AXI_RM_BCM00_CK_AND `i_axi_DW_AXI_RM_BCM00_CK_AND
`endif 

`ifdef i_axi_DW_AXI_RM_BCM00_CK_BUF
  `define DW_AXI_RM_BCM00_CK_BUF `i_axi_DW_AXI_RM_BCM00_CK_BUF
`endif 

`ifdef i_axi_DW_AXI_RM_BCM00_CK_GT_LAT
  `define DW_AXI_RM_BCM00_CK_GT_LAT `i_axi_DW_AXI_RM_BCM00_CK_GT_LAT
`endif 

`ifdef i_axi_DW_AXI_RM_BCM00_CK_MX
  `define DW_AXI_RM_BCM00_CK_MX `i_axi_DW_AXI_RM_BCM00_CK_MX
`endif 

`ifdef i_axi_DW_AXI_RM_BCM00_CK_OR
  `define DW_AXI_RM_BCM00_CK_OR `i_axi_DW_AXI_RM_BCM00_CK_OR
`endif 

`ifdef i_axi_DW_AXI_RM_BCM00_MAJ
  `define DW_AXI_RM_BCM00_MAJ `i_axi_DW_AXI_RM_BCM00_MAJ
`endif 

`ifdef i_axi_DW_AXI_RM_BCM00_MX
  `define DW_AXI_RM_BCM00_MX `i_axi_DW_AXI_RM_BCM00_MX
`endif 

`ifdef i_axi_DW_AXI_RM_BCM00_OR
  `define DW_AXI_RM_BCM00_OR `i_axi_DW_AXI_RM_BCM00_OR
`endif 

`ifdef i_axi_DW_AXI_RM_BCM01
  `define DW_AXI_RM_BCM01 `i_axi_DW_AXI_RM_BCM01
`endif 

`ifdef i_axi_DW_AXI_RM_BCM02
  `define DW_AXI_RM_BCM02 `i_axi_DW_AXI_RM_BCM02
`endif 

`ifdef i_axi_DW_AXI_RM_BCM03
  `define DW_AXI_RM_BCM03 `i_axi_DW_AXI_RM_BCM03
`endif 

`ifdef i_axi_DW_AXI_RM_BCM04
  `define DW_AXI_RM_BCM04 `i_axi_DW_AXI_RM_BCM04
`endif 

`ifdef i_axi_DW_AXI_RM_BCM05
  `define DW_AXI_RM_BCM05 `i_axi_DW_AXI_RM_BCM05
`endif 

`ifdef i_axi_DW_AXI_RM_BCM05_ATV
  `define DW_AXI_RM_BCM05_ATV `i_axi_DW_AXI_RM_BCM05_ATV
`endif 

`ifdef i_axi_DW_AXI_RM_BCM05_CF
  `define DW_AXI_RM_BCM05_CF `i_axi_DW_AXI_RM_BCM05_CF
`endif 

`ifdef i_axi_DW_AXI_RM_BCM05_EF
  `define DW_AXI_RM_BCM05_EF `i_axi_DW_AXI_RM_BCM05_EF
`endif 

`ifdef i_axi_DW_AXI_RM_BCM05_EF_ATV
  `define DW_AXI_RM_BCM05_EF_ATV `i_axi_DW_AXI_RM_BCM05_EF_ATV
`endif 

`ifdef i_axi_DW_AXI_RM_BCM06
  `define DW_AXI_RM_BCM06 `i_axi_DW_AXI_RM_BCM06
`endif 

`ifdef i_axi_DW_AXI_RM_BCM06_ATV
  `define DW_AXI_RM_BCM06_ATV `i_axi_DW_AXI_RM_BCM06_ATV
`endif 

`ifdef i_axi_DW_AXI_RM_BCM07
  `define DW_AXI_RM_BCM07 `i_axi_DW_AXI_RM_BCM07
`endif 

`ifdef i_axi_DW_AXI_RM_BCM07_ATV
  `define DW_AXI_RM_BCM07_ATV `i_axi_DW_AXI_RM_BCM07_ATV
`endif 

`ifdef i_axi_DW_AXI_RM_BCM07_EF
  `define DW_AXI_RM_BCM07_EF `i_axi_DW_AXI_RM_BCM07_EF
`endif 

`ifdef i_axi_DW_AXI_RM_BCM07_EF_ATV
  `define DW_AXI_RM_BCM07_EF_ATV `i_axi_DW_AXI_RM_BCM07_EF_ATV
`endif 

`ifdef i_axi_DW_AXI_RM_BCM07_EFES
  `define DW_AXI_RM_BCM07_EFES `i_axi_DW_AXI_RM_BCM07_EFES
`endif 

`ifdef i_axi_DW_AXI_RM_BCM07_RS
  `define DW_AXI_RM_BCM07_RS `i_axi_DW_AXI_RM_BCM07_RS
`endif 

`ifdef i_axi_DW_AXI_RM_BCM08
  `define DW_AXI_RM_BCM08 `i_axi_DW_AXI_RM_BCM08
`endif 

`ifdef i_axi_DW_AXI_RM_BCM09
  `define DW_AXI_RM_BCM09 `i_axi_DW_AXI_RM_BCM09
`endif 

`ifdef i_axi_DW_AXI_RM_BCM09_DP
  `define DW_AXI_RM_BCM09_DP `i_axi_DW_AXI_RM_BCM09_DP
`endif 

`ifdef i_axi_DW_AXI_RM_BCM09_ECC
  `define DW_AXI_RM_BCM09_ECC `i_axi_DW_AXI_RM_BCM09_ECC
`endif 

`ifdef i_axi_DW_AXI_RM_BCM10
  `define DW_AXI_RM_BCM10 `i_axi_DW_AXI_RM_BCM10
`endif 

`ifdef i_axi_DW_AXI_RM_BCM11
  `define DW_AXI_RM_BCM11 `i_axi_DW_AXI_RM_BCM11
`endif 

`ifdef i_axi_DW_AXI_RM_BCM12
  `define DW_AXI_RM_BCM12 `i_axi_DW_AXI_RM_BCM12
`endif 

`ifdef i_axi_DW_AXI_RM_BCM14
  `define DW_AXI_RM_BCM14 `i_axi_DW_AXI_RM_BCM14
`endif 

`ifdef i_axi_DW_AXI_RM_BCM15
  `define DW_AXI_RM_BCM15 `i_axi_DW_AXI_RM_BCM15
`endif 

`ifdef i_axi_DW_AXI_RM_BCM16
  `define DW_AXI_RM_BCM16 `i_axi_DW_AXI_RM_BCM16
`endif 

`ifdef i_axi_DW_AXI_RM_BCM17
  `define DW_AXI_RM_BCM17 `i_axi_DW_AXI_RM_BCM17
`endif 

`ifdef i_axi_DW_AXI_RM_BCM18_GEN
  `define DW_AXI_RM_BCM18_GEN `i_axi_DW_AXI_RM_BCM18_GEN
`endif 

`ifdef i_axi_DW_AXI_RM_BCM18_MON
  `define DW_AXI_RM_BCM18_MON `i_axi_DW_AXI_RM_BCM18_MON
`endif 

`ifdef i_axi_DW_AXI_RM_BCM18_PGEN
  `define DW_AXI_RM_BCM18_PGEN `i_axi_DW_AXI_RM_BCM18_PGEN
`endif 

`ifdef i_axi_DW_AXI_RM_BCM18_PGENA
  `define DW_AXI_RM_BCM18_PGENA `i_axi_DW_AXI_RM_BCM18_PGENA
`endif 

`ifdef i_axi_DW_AXI_RM_BCM18_PMON
  `define DW_AXI_RM_BCM18_PMON `i_axi_DW_AXI_RM_BCM18_PMON
`endif 

`ifdef i_axi_DW_AXI_RM_BCM18_RS
  `define DW_AXI_RM_BCM18_RS `i_axi_DW_AXI_RM_BCM18_RS
`endif 

`ifdef i_axi_DW_AXI_RM_BCM19_INTR
  `define DW_AXI_RM_BCM19_INTR `i_axi_DW_AXI_RM_BCM19_INTR
`endif 

`ifdef i_axi_DW_AXI_RM_BCM19_TRGT
  `define DW_AXI_RM_BCM19_TRGT `i_axi_DW_AXI_RM_BCM19_TRGT
`endif 

`ifdef i_axi_DW_AXI_RM_BCM21
  `define DW_AXI_RM_BCM21 `i_axi_DW_AXI_RM_BCM21
`endif 

`ifdef i_axi_DW_AXI_RM_BCM21_ATV
  `define DW_AXI_RM_BCM21_ATV `i_axi_DW_AXI_RM_BCM21_ATV
`endif 

`ifdef i_axi_DW_AXI_RM_BCM21_NEO
  `define DW_AXI_RM_BCM21_NEO `i_axi_DW_AXI_RM_BCM21_NEO
`endif 

`ifdef i_axi_DW_AXI_RM_BCM21_TGL
  `define DW_AXI_RM_BCM21_TGL `i_axi_DW_AXI_RM_BCM21_TGL
`endif 

`ifdef i_axi_DW_AXI_RM_BCM22
  `define DW_AXI_RM_BCM22 `i_axi_DW_AXI_RM_BCM22
`endif 

`ifdef i_axi_DW_AXI_RM_BCM22_ATV
  `define DW_AXI_RM_BCM22_ATV `i_axi_DW_AXI_RM_BCM22_ATV
`endif 

`ifdef i_axi_DW_AXI_RM_BCM23
  `define DW_AXI_RM_BCM23 `i_axi_DW_AXI_RM_BCM23
`endif 

`ifdef i_axi_DW_AXI_RM_BCM23_ATV
  `define DW_AXI_RM_BCM23_ATV `i_axi_DW_AXI_RM_BCM23_ATV
`endif 

`ifdef i_axi_DW_AXI_RM_BCM23_C
  `define DW_AXI_RM_BCM23_C `i_axi_DW_AXI_RM_BCM23_C
`endif 

`ifdef i_axi_DW_AXI_RM_BCM24
  `define DW_AXI_RM_BCM24 `i_axi_DW_AXI_RM_BCM24
`endif 

`ifdef i_axi_DW_AXI_RM_BCM24_AP
  `define DW_AXI_RM_BCM24_AP `i_axi_DW_AXI_RM_BCM24_AP
`endif 

`ifdef i_axi_DW_AXI_RM_BCM25
  `define DW_AXI_RM_BCM25 `i_axi_DW_AXI_RM_BCM25
`endif 

`ifdef i_axi_DW_AXI_RM_BCM25_ATV
  `define DW_AXI_RM_BCM25_ATV `i_axi_DW_AXI_RM_BCM25_ATV
`endif 

`ifdef i_axi_DW_AXI_RM_BCM25_C
  `define DW_AXI_RM_BCM25_C `i_axi_DW_AXI_RM_BCM25_C
`endif 

`ifdef i_axi_DW_AXI_RM_BCM26
  `define DW_AXI_RM_BCM26 `i_axi_DW_AXI_RM_BCM26
`endif 

`ifdef i_axi_DW_AXI_RM_BCM26_ATV
  `define DW_AXI_RM_BCM26_ATV `i_axi_DW_AXI_RM_BCM26_ATV
`endif 

`ifdef i_axi_DW_AXI_RM_BCM27
  `define DW_AXI_RM_BCM27 `i_axi_DW_AXI_RM_BCM27
`endif 

`ifdef i_axi_DW_AXI_RM_BCM28
  `define DW_AXI_RM_BCM28 `i_axi_DW_AXI_RM_BCM28
`endif 

`ifdef i_axi_DW_AXI_RM_BCM29
  `define DW_AXI_RM_BCM29 `i_axi_DW_AXI_RM_BCM29
`endif 

`ifdef i_axi_DW_AXI_RM_BCM31_P2D_FIFOMEM
  `define DW_AXI_RM_BCM31_P2D_FIFOMEM `i_axi_DW_AXI_RM_BCM31_P2D_FIFOMEM
`endif 

`ifdef i_axi_DW_AXI_RM_BCM31_P2D_RD
  `define DW_AXI_RM_BCM31_P2D_RD `i_axi_DW_AXI_RM_BCM31_P2D_RD
`endif 

`ifdef i_axi_DW_AXI_RM_BCM31_P2D_WR
  `define DW_AXI_RM_BCM31_P2D_WR `i_axi_DW_AXI_RM_BCM31_P2D_WR
`endif 

`ifdef i_axi_DW_AXI_RM_BCM32_A
  `define DW_AXI_RM_BCM32_A `i_axi_DW_AXI_RM_BCM32_A
`endif 

`ifdef i_axi_DW_AXI_RM_BCM32_C
  `define DW_AXI_RM_BCM32_C `i_axi_DW_AXI_RM_BCM32_C
`endif 

`ifdef i_axi_DW_AXI_RM_BCM33_63_7_64_0
  `define DW_AXI_RM_BCM33_63_7_64_0 `i_axi_DW_AXI_RM_BCM33_63_7_64_0
`endif 

`ifdef i_axi_DW_AXI_RM_BCM35
  `define DW_AXI_RM_BCM35 `i_axi_DW_AXI_RM_BCM35
`endif 

`ifdef i_axi_DW_AXI_RM_BCM35_T
  `define DW_AXI_RM_BCM35_T `i_axi_DW_AXI_RM_BCM35_T
`endif 

`ifdef i_axi_DW_AXI_RM_BCM36
  `define DW_AXI_RM_BCM36 `i_axi_DW_AXI_RM_BCM36
`endif 

`ifdef i_axi_DW_AXI_RM_BCM36_ACK
  `define DW_AXI_RM_BCM36_ACK `i_axi_DW_AXI_RM_BCM36_ACK
`endif 

`ifdef i_axi_DW_AXI_RM_BCM36_NHS
  `define DW_AXI_RM_BCM36_NHS `i_axi_DW_AXI_RM_BCM36_NHS
`endif 

`ifdef i_axi_DW_AXI_RM_BCM36_TGL
  `define DW_AXI_RM_BCM36_TGL `i_axi_DW_AXI_RM_BCM36_TGL
`endif 

`ifdef i_axi_DW_AXI_RM_BCM36_TGL_DO
  `define DW_AXI_RM_BCM36_TGL_DO `i_axi_DW_AXI_RM_BCM36_TGL_DO
`endif 

`ifdef i_axi_DW_AXI_RM_BCM36_TGL_PLS
  `define DW_AXI_RM_BCM36_TGL_PLS `i_axi_DW_AXI_RM_BCM36_TGL_PLS
`endif 

`ifdef i_axi_DW_AXI_RM_BCM36_TGL_PLS_DO
  `define DW_AXI_RM_BCM36_TGL_PLS_DO `i_axi_DW_AXI_RM_BCM36_TGL_PLS_DO
`endif 

`ifdef i_axi_DW_AXI_RM_BCM37
  `define DW_AXI_RM_BCM37 `i_axi_DW_AXI_RM_BCM37
`endif 

`ifdef i_axi_DW_AXI_RM_BCM38
  `define DW_AXI_RM_BCM38 `i_axi_DW_AXI_RM_BCM38
`endif 

`ifdef i_axi_DW_AXI_RM_BCM38_ADP
  `define DW_AXI_RM_BCM38_ADP `i_axi_DW_AXI_RM_BCM38_ADP
`endif 

`ifdef i_axi_DW_AXI_RM_BCM38_AP
  `define DW_AXI_RM_BCM38_AP `i_axi_DW_AXI_RM_BCM38_AP
`endif 

`ifdef i_axi_DW_AXI_RM_BCM38_ECC
  `define DW_AXI_RM_BCM38_ECC `i_axi_DW_AXI_RM_BCM38_ECC
`endif 

`ifdef i_axi_DW_AXI_RM_BCM39
  `define DW_AXI_RM_BCM39 `i_axi_DW_AXI_RM_BCM39
`endif 

`ifdef i_axi_DW_AXI_RM_BCM40
  `define DW_AXI_RM_BCM40 `i_axi_DW_AXI_RM_BCM40
`endif 

`ifdef i_axi_DW_AXI_RM_BCM41
  `define DW_AXI_RM_BCM41 `i_axi_DW_AXI_RM_BCM41
`endif 

`ifdef i_axi_DW_AXI_RM_BCM41_NEO
  `define DW_AXI_RM_BCM41_NEO `i_axi_DW_AXI_RM_BCM41_NEO
`endif 

`ifdef i_axi_DW_AXI_RM_BCM43
  `define DW_AXI_RM_BCM43 `i_axi_DW_AXI_RM_BCM43
`endif 

`ifdef i_axi_DW_AXI_RM_BCM43_NRO
  `define DW_AXI_RM_BCM43_NRO `i_axi_DW_AXI_RM_BCM43_NRO
`endif 

`ifdef i_axi_DW_AXI_RM_BCM44
  `define DW_AXI_RM_BCM44 `i_axi_DW_AXI_RM_BCM44
`endif 

`ifdef i_axi_DW_AXI_RM_BCM44_NRO
  `define DW_AXI_RM_BCM44_NRO `i_axi_DW_AXI_RM_BCM44_NRO
`endif 

`ifdef i_axi_DW_AXI_RM_BCM45_GN_D_A
  `define DW_AXI_RM_BCM45_GN_D_A `i_axi_DW_AXI_RM_BCM45_GN_D_A
`endif 

`ifdef i_axi_DW_AXI_RM_BCM45_GN_D_AA
  `define DW_AXI_RM_BCM45_GN_D_AA `i_axi_DW_AXI_RM_BCM45_GN_D_AA
`endif 

`ifdef i_axi_DW_AXI_RM_BCM45_GN_D_B
  `define DW_AXI_RM_BCM45_GN_D_B `i_axi_DW_AXI_RM_BCM45_GN_D_B
`endif 

`ifdef i_axi_DW_AXI_RM_BCM45_GN_D_C
  `define DW_AXI_RM_BCM45_GN_D_C `i_axi_DW_AXI_RM_BCM45_GN_D_C
`endif 

`ifdef i_axi_DW_AXI_RM_BCM45_GN_D_D
  `define DW_AXI_RM_BCM45_GN_D_D `i_axi_DW_AXI_RM_BCM45_GN_D_D
`endif 

`ifdef i_axi_DW_AXI_RM_BCM45_GN_D_E
  `define DW_AXI_RM_BCM45_GN_D_E `i_axi_DW_AXI_RM_BCM45_GN_D_E
`endif 

`ifdef i_axi_DW_AXI_RM_BCM45_GN_D_F
  `define DW_AXI_RM_BCM45_GN_D_F `i_axi_DW_AXI_RM_BCM45_GN_D_F
`endif 

`ifdef i_axi_DW_AXI_RM_BCM45_MN_D_A
  `define DW_AXI_RM_BCM45_MN_D_A `i_axi_DW_AXI_RM_BCM45_MN_D_A
`endif 

`ifdef i_axi_DW_AXI_RM_BCM45_MN_D_AA
  `define DW_AXI_RM_BCM45_MN_D_AA `i_axi_DW_AXI_RM_BCM45_MN_D_AA
`endif 

`ifdef i_axi_DW_AXI_RM_BCM45_MN_D_B
  `define DW_AXI_RM_BCM45_MN_D_B `i_axi_DW_AXI_RM_BCM45_MN_D_B
`endif 

`ifdef i_axi_DW_AXI_RM_BCM45_MN_D_C
  `define DW_AXI_RM_BCM45_MN_D_C `i_axi_DW_AXI_RM_BCM45_MN_D_C
`endif 

`ifdef i_axi_DW_AXI_RM_BCM45_MN_D_D
  `define DW_AXI_RM_BCM45_MN_D_D `i_axi_DW_AXI_RM_BCM45_MN_D_D
`endif 

`ifdef i_axi_DW_AXI_RM_BCM45_MN_D_E
  `define DW_AXI_RM_BCM45_MN_D_E `i_axi_DW_AXI_RM_BCM45_MN_D_E
`endif 

`ifdef i_axi_DW_AXI_RM_BCM45_MN_D_F
  `define DW_AXI_RM_BCM45_MN_D_F `i_axi_DW_AXI_RM_BCM45_MN_D_F
`endif 

`ifdef i_axi_DW_AXI_RM_BCM46_A
  `define DW_AXI_RM_BCM46_A `i_axi_DW_AXI_RM_BCM46_A
`endif 

`ifdef i_axi_DW_AXI_RM_BCM46_AA
  `define DW_AXI_RM_BCM46_AA `i_axi_DW_AXI_RM_BCM46_AA
`endif 

`ifdef i_axi_DW_AXI_RM_BCM46_B
  `define DW_AXI_RM_BCM46_B `i_axi_DW_AXI_RM_BCM46_B
`endif 

`ifdef i_axi_DW_AXI_RM_BCM46_B_32A
  `define DW_AXI_RM_BCM46_B_32A `i_axi_DW_AXI_RM_BCM46_B_32A
`endif 

`ifdef i_axi_DW_AXI_RM_BCM46_C
  `define DW_AXI_RM_BCM46_C `i_axi_DW_AXI_RM_BCM46_C
`endif 

`ifdef i_axi_DW_AXI_RM_BCM46_C_64A
  `define DW_AXI_RM_BCM46_C_64A `i_axi_DW_AXI_RM_BCM46_C_64A
`endif 

`ifdef i_axi_DW_AXI_RM_BCM46_D
  `define DW_AXI_RM_BCM46_D `i_axi_DW_AXI_RM_BCM46_D
`endif 

`ifdef i_axi_DW_AXI_RM_BCM46_D_128A
  `define DW_AXI_RM_BCM46_D_128A `i_axi_DW_AXI_RM_BCM46_D_128A
`endif 

`ifdef i_axi_DW_AXI_RM_BCM46_E
  `define DW_AXI_RM_BCM46_E `i_axi_DW_AXI_RM_BCM46_E
`endif 

`ifdef i_axi_DW_AXI_RM_BCM46_F
  `define DW_AXI_RM_BCM46_F `i_axi_DW_AXI_RM_BCM46_F
`endif 

`ifdef i_axi_DW_AXI_RM_BCM46_X
  `define DW_AXI_RM_BCM46_X `i_axi_DW_AXI_RM_BCM46_X
`endif 

`ifdef i_axi_DW_AXI_RM_BCM47
  `define DW_AXI_RM_BCM47 `i_axi_DW_AXI_RM_BCM47
`endif 

`ifdef i_axi_DW_AXI_RM_BCM48
  `define DW_AXI_RM_BCM48 `i_axi_DW_AXI_RM_BCM48
`endif 

`ifdef i_axi_DW_AXI_RM_BCM48_DM
  `define DW_AXI_RM_BCM48_DM `i_axi_DW_AXI_RM_BCM48_DM
`endif 

`ifdef i_axi_DW_AXI_RM_BCM48_SV
  `define DW_AXI_RM_BCM48_SV `i_axi_DW_AXI_RM_BCM48_SV
`endif 

`ifdef i_axi_DW_AXI_RM_BCM49
  `define DW_AXI_RM_BCM49 `i_axi_DW_AXI_RM_BCM49
`endif 

`ifdef i_axi_DW_AXI_RM_BCM49_SV
  `define DW_AXI_RM_BCM49_SV `i_axi_DW_AXI_RM_BCM49_SV
`endif 

`ifdef i_axi_DW_AXI_RM_BCM50
  `define DW_AXI_RM_BCM50 `i_axi_DW_AXI_RM_BCM50
`endif 

`ifdef i_axi_DW_AXI_RM_BCM51
  `define DW_AXI_RM_BCM51 `i_axi_DW_AXI_RM_BCM51
`endif 

`ifdef i_axi_DW_AXI_RM_BCM52
  `define DW_AXI_RM_BCM52 `i_axi_DW_AXI_RM_BCM52
`endif 

`ifdef i_axi_DW_AXI_RM_BCM53
  `define DW_AXI_RM_BCM53 `i_axi_DW_AXI_RM_BCM53
`endif 

`ifdef i_axi_DW_AXI_RM_BCM54
  `define DW_AXI_RM_BCM54 `i_axi_DW_AXI_RM_BCM54
`endif 

`ifdef i_axi_DW_AXI_RM_BCM55
  `define DW_AXI_RM_BCM55 `i_axi_DW_AXI_RM_BCM55
`endif 

`ifdef i_axi_DW_AXI_RM_BCM55_C
  `define DW_AXI_RM_BCM55_C `i_axi_DW_AXI_RM_BCM55_C
`endif 

`ifdef i_axi_DW_AXI_RM_BCM56
  `define DW_AXI_RM_BCM56 `i_axi_DW_AXI_RM_BCM56
`endif 

`ifdef i_axi_DW_AXI_RM_BCM57
  `define DW_AXI_RM_BCM57 `i_axi_DW_AXI_RM_BCM57
`endif 

`ifdef i_axi_DW_AXI_RM_BCM57_ATV
  `define DW_AXI_RM_BCM57_ATV `i_axi_DW_AXI_RM_BCM57_ATV
`endif 

`ifdef i_axi_DW_AXI_RM_BCM58
  `define DW_AXI_RM_BCM58 `i_axi_DW_AXI_RM_BCM58
`endif 

`ifdef i_axi_DW_AXI_RM_BCM58_ATV
  `define DW_AXI_RM_BCM58_ATV `i_axi_DW_AXI_RM_BCM58_ATV
`endif 

`ifdef i_axi_DW_AXI_RM_BCM59
  `define DW_AXI_RM_BCM59 `i_axi_DW_AXI_RM_BCM59
`endif 

`ifdef i_axi_DW_AXI_RM_BCM60
  `define DW_AXI_RM_BCM60 `i_axi_DW_AXI_RM_BCM60
`endif 

`ifdef i_axi_DW_AXI_RM_BCM62
  `define DW_AXI_RM_BCM62 `i_axi_DW_AXI_RM_BCM62
`endif 

`ifdef i_axi_DW_AXI_RM_BCM63
  `define DW_AXI_RM_BCM63 `i_axi_DW_AXI_RM_BCM63
`endif 

`ifdef i_axi_DW_AXI_RM_BCM64
  `define DW_AXI_RM_BCM64 `i_axi_DW_AXI_RM_BCM64
`endif 

`ifdef i_axi_DW_AXI_RM_BCM64_TD
  `define DW_AXI_RM_BCM64_TD `i_axi_DW_AXI_RM_BCM64_TD
`endif 

`ifdef i_axi_DW_AXI_RM_BCM65
  `define DW_AXI_RM_BCM65 `i_axi_DW_AXI_RM_BCM65
`endif 

`ifdef i_axi_DW_AXI_RM_BCM65_ATV
  `define DW_AXI_RM_BCM65_ATV `i_axi_DW_AXI_RM_BCM65_ATV
`endif 

`ifdef i_axi_DW_AXI_RM_BCM65_TD
  `define DW_AXI_RM_BCM65_TD `i_axi_DW_AXI_RM_BCM65_TD
`endif 

`ifdef i_axi_DW_AXI_RM_BCM66
  `define DW_AXI_RM_BCM66 `i_axi_DW_AXI_RM_BCM66
`endif 

`ifdef i_axi_DW_AXI_RM_BCM66_ATV
  `define DW_AXI_RM_BCM66_ATV `i_axi_DW_AXI_RM_BCM66_ATV
`endif 

`ifdef i_axi_DW_AXI_RM_BCM66_DMS
  `define DW_AXI_RM_BCM66_DMS `i_axi_DW_AXI_RM_BCM66_DMS
`endif 

`ifdef i_axi_DW_AXI_RM_BCM66_DMS_ATV
  `define DW_AXI_RM_BCM66_DMS_ATV `i_axi_DW_AXI_RM_BCM66_DMS_ATV
`endif 

`ifdef i_axi_DW_AXI_RM_BCM66_EFES
  `define DW_AXI_RM_BCM66_EFES `i_axi_DW_AXI_RM_BCM66_EFES
`endif 

`ifdef i_axi_DW_AXI_RM_BCM66_PR
  `define DW_AXI_RM_BCM66_PR `i_axi_DW_AXI_RM_BCM66_PR
`endif 

`ifdef i_axi_DW_AXI_RM_BCM66_WAE
  `define DW_AXI_RM_BCM66_WAE `i_axi_DW_AXI_RM_BCM66_WAE
`endif 

`ifdef i_axi_DW_AXI_RM_BCM66_WAE_ATV
  `define DW_AXI_RM_BCM66_WAE_ATV `i_axi_DW_AXI_RM_BCM66_WAE_ATV
`endif 

`ifdef i_axi_DW_AXI_RM_BCM68_63_7_0
  `define DW_AXI_RM_BCM68_63_7_0 `i_axi_DW_AXI_RM_BCM68_63_7_0
`endif 

`ifdef i_axi_DW_AXI_RM_BCM69_63_7_0
  `define DW_AXI_RM_BCM69_63_7_0 `i_axi_DW_AXI_RM_BCM69_63_7_0
`endif 

`ifdef i_axi_DW_AXI_RM_BCM70_63_7_0_0
  `define DW_AXI_RM_BCM70_63_7_0_0 `i_axi_DW_AXI_RM_BCM70_63_7_0_0
`endif 

`ifdef i_axi_DW_AXI_RM_BCM71
  `define DW_AXI_RM_BCM71 `i_axi_DW_AXI_RM_BCM71
`endif 

`ifdef i_axi_DW_AXI_RM_BCM72
  `define DW_AXI_RM_BCM72 `i_axi_DW_AXI_RM_BCM72
`endif 

`ifdef i_axi_DW_AXI_RM_BCM74
  `define DW_AXI_RM_BCM74 `i_axi_DW_AXI_RM_BCM74
`endif 

`ifdef i_axi_DW_AXI_RM_BCM76
  `define DW_AXI_RM_BCM76 `i_axi_DW_AXI_RM_BCM76
`endif 

`ifdef i_axi_DW_AXI_RM_BCM77
  `define DW_AXI_RM_BCM77 `i_axi_DW_AXI_RM_BCM77
`endif 

`ifdef i_axi_DW_AXI_RM_BCM78
  `define DW_AXI_RM_BCM78 `i_axi_DW_AXI_RM_BCM78
`endif 

`ifdef i_axi_DW_AXI_RM_BCM79
  `define DW_AXI_RM_BCM79 `i_axi_DW_AXI_RM_BCM79
`endif 

`ifdef i_axi_DW_AXI_RM_BCM79_MO
  `define DW_AXI_RM_BCM79_MO `i_axi_DW_AXI_RM_BCM79_MO
`endif 

`ifdef i_axi_DW_AXI_RM_BCM83_GEN
  `define DW_AXI_RM_BCM83_GEN `i_axi_DW_AXI_RM_BCM83_GEN
`endif 

`ifdef i_axi_DW_AXI_RM_BCM84_MON
  `define DW_AXI_RM_BCM84_MON `i_axi_DW_AXI_RM_BCM84_MON
`endif 

`ifdef i_axi_DW_AXI_RM_BCM85
  `define DW_AXI_RM_BCM85 `i_axi_DW_AXI_RM_BCM85
`endif 

`ifdef i_axi_DW_AXI_RM_BCM86
  `define DW_AXI_RM_BCM86 `i_axi_DW_AXI_RM_BCM86
`endif 

`ifdef i_axi_DW_AXI_RM_BCM87
  `define DW_AXI_RM_BCM87 `i_axi_DW_AXI_RM_BCM87
`endif 

`ifdef i_axi_DW_AXI_RM_BCM90
  `define DW_AXI_RM_BCM90 `i_axi_DW_AXI_RM_BCM90
`endif 

`ifdef i_axi_DW_AXI_RM_BCM91
  `define DW_AXI_RM_BCM91 `i_axi_DW_AXI_RM_BCM91
`endif 

`ifdef i_axi_DW_AXI_RM_BCM92
  `define DW_AXI_RM_BCM92 `i_axi_DW_AXI_RM_BCM92
`endif 

`ifdef i_axi_DW_AXI_RM_BCM92_AD
  `define DW_AXI_RM_BCM92_AD `i_axi_DW_AXI_RM_BCM92_AD
`endif 

`ifdef i_axi_DW_AXI_RM_BCM92_AD_DO
  `define DW_AXI_RM_BCM92_AD_DO `i_axi_DW_AXI_RM_BCM92_AD_DO
`endif 

`ifdef i_axi_DW_AXI_RM_BCM92_RD
  `define DW_AXI_RM_BCM92_RD `i_axi_DW_AXI_RM_BCM92_RD
`endif 

`ifdef i_axi_DW_AXI_RM_BCM92_RD_AD
  `define DW_AXI_RM_BCM92_RD_AD `i_axi_DW_AXI_RM_BCM92_RD_AD
`endif 

`ifdef i_axi_DW_AXI_RM_BCM92_RD_AD_DO
  `define DW_AXI_RM_BCM92_RD_AD_DO `i_axi_DW_AXI_RM_BCM92_RD_AD_DO
`endif 

`ifdef i_axi_DW_AXI_RM_BCM92_RD_DO
  `define DW_AXI_RM_BCM92_RD_DO `i_axi_DW_AXI_RM_BCM92_RD_DO
`endif 

`ifdef i_axi_DW_AXI_RM_BCM93
  `define DW_AXI_RM_BCM93 `i_axi_DW_AXI_RM_BCM93
`endif 

`ifdef i_axi_DW_AXI_RM_BCM93_NDSVA
  `define DW_AXI_RM_BCM93_NDSVA `i_axi_DW_AXI_RM_BCM93_NDSVA
`endif 

`ifdef i_axi_DW_AXI_RM_BCM94
  `define DW_AXI_RM_BCM94 `i_axi_DW_AXI_RM_BCM94
`endif 

`ifdef i_axi_DW_AXI_RM_BCM95
  `define DW_AXI_RM_BCM95 `i_axi_DW_AXI_RM_BCM95
`endif 

`ifdef i_axi_DW_AXI_RM_BCM95_E
  `define DW_AXI_RM_BCM95_E `i_axi_DW_AXI_RM_BCM95_E
`endif 

`ifdef i_axi_DW_AXI_RM_BCM95_I
  `define DW_AXI_RM_BCM95_I `i_axi_DW_AXI_RM_BCM95_I
`endif 

`ifdef i_axi_DW_AXI_RM_BCM95_IE
  `define DW_AXI_RM_BCM95_IE `i_axi_DW_AXI_RM_BCM95_IE
`endif 

`ifdef i_axi_DW_AXI_RM_BCM95_NE
  `define DW_AXI_RM_BCM95_NE `i_axi_DW_AXI_RM_BCM95_NE
`endif 

`ifdef i_axi_DW_AXI_RM_BCM95_NE_E
  `define DW_AXI_RM_BCM95_NE_E `i_axi_DW_AXI_RM_BCM95_NE_E
`endif 

`ifdef i_axi_DW_AXI_RM_BCM95_NE_I
  `define DW_AXI_RM_BCM95_NE_I `i_axi_DW_AXI_RM_BCM95_NE_I
`endif 

`ifdef i_axi_DW_AXI_RM_BCM95_NE_IE
  `define DW_AXI_RM_BCM95_NE_IE `i_axi_DW_AXI_RM_BCM95_NE_IE
`endif 

`ifdef i_axi_DW_AXI_RM_BCM98
  `define DW_AXI_RM_BCM98 `i_axi_DW_AXI_RM_BCM98
`endif 

`ifdef i_axi_DW_AXI_RM_BCM99
  `define DW_AXI_RM_BCM99 `i_axi_DW_AXI_RM_BCM99
`endif 

`ifdef i_axi_DW_AXI_RM_BCM99_3
  `define DW_AXI_RM_BCM99_3 `i_axi_DW_AXI_RM_BCM99_3
`endif 

`ifdef i_axi_DW_AXI_RM_BCM99_4
  `define DW_AXI_RM_BCM99_4 `i_axi_DW_AXI_RM_BCM99_4
`endif 

`ifdef i_axi_DW_AXI_RM_BCM99_N
  `define DW_AXI_RM_BCM99_N `i_axi_DW_AXI_RM_BCM99_N
`endif 

`ifdef i_axi_DW_AXI_RM_BVM01
  `define DW_AXI_RM_BVM01 `i_axi_DW_AXI_RM_BVM01
`endif 

`ifdef i_axi_DW_AXI_RM_BVM02
  `define DW_AXI_RM_BVM02 `i_axi_DW_AXI_RM_BVM02
`endif 

`ifdef i_axi_DW_AXI_RM_SVA01
  `define DW_AXI_RM_SVA01 `i_axi_DW_AXI_RM_SVA01
`endif 

`ifdef i_axi_DW_AXI_RM_SVA02
  `define DW_AXI_RM_SVA02 `i_axi_DW_AXI_RM_SVA02
`endif 

`ifdef i_axi_DW_AXI_RM_SVA03
  `define DW_AXI_RM_SVA03 `i_axi_DW_AXI_RM_SVA03
`endif 

`ifdef i_axi_DW_AXI_RM_SVA04
  `define DW_AXI_RM_SVA04 `i_axi_DW_AXI_RM_SVA04
`endif 

`ifdef i_axi_DW_AXI_RM_SVA05
  `define DW_AXI_RM_SVA05 `i_axi_DW_AXI_RM_SVA05
`endif 

`ifdef i_axi_DW_AXI_RM_SVA06
  `define DW_AXI_RM_SVA06 `i_axi_DW_AXI_RM_SVA06
`endif 

`ifdef i_axi_DW_AXI_RM_SVA07
  `define DW_AXI_RM_SVA07 `i_axi_DW_AXI_RM_SVA07
`endif 

`ifdef i_axi_DW_AXI_RM_SVA08
  `define DW_AXI_RM_SVA08 `i_axi_DW_AXI_RM_SVA08
`endif 

`ifdef i_axi_DW_AXI_RM_SVA09
  `define DW_AXI_RM_SVA09 `i_axi_DW_AXI_RM_SVA09
`endif 

`ifdef i_axi_DW_AXI_RM_SVA10
  `define DW_AXI_RM_SVA10 `i_axi_DW_AXI_RM_SVA10
`endif 

`ifdef i_axi_DW_AXI_RM_SVA11
  `define DW_AXI_RM_SVA11 `i_axi_DW_AXI_RM_SVA11
`endif 

`ifdef i_axi_DW_AXI_RM_SVA12_A
  `define DW_AXI_RM_SVA12_A `i_axi_DW_AXI_RM_SVA12_A
`endif 

`ifdef i_axi_DW_AXI_RM_SVA12_B
  `define DW_AXI_RM_SVA12_B `i_axi_DW_AXI_RM_SVA12_B
`endif 

`ifdef i_axi_DW_AXI_RM_SVA12_C
  `define DW_AXI_RM_SVA12_C `i_axi_DW_AXI_RM_SVA12_C
`endif 

`ifdef i_axi_DW_AXI_RM_SVA99
  `define DW_AXI_RM_SVA99 `i_axi_DW_AXI_RM_SVA99
`endif 

`ifdef i_axi___GUARD__DW_AXI_ALL_INCLUDES__VH__
  `define __GUARD__DW_AXI_ALL_INCLUDES__VH__ `i_axi___GUARD__DW_AXI_ALL_INCLUDES__VH__
`endif 

`ifdef i_axi_DW_HOLD_MUX_DELAY
  `define DW_HOLD_MUX_DELAY `i_axi_DW_HOLD_MUX_DELAY
`endif 

`ifdef i_axi_DW_SETUP_MUX_DELAY
  `define DW_SETUP_MUX_DELAY `i_axi_DW_SETUP_MUX_DELAY
`endif 

`ifdef i_axi_cb_dummy_parameter_definition
  `define cb_dummy_parameter_definition `i_axi_cb_dummy_parameter_definition
`endif 

