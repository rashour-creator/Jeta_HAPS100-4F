`define __GUARD__DW_AXI_CC_CONSTANTS__VH__
`define AXI_USE_RANDOM_SEED 0
`define AXI_SEED 32'h1
`define USE_FOUNDATION 1
`define AXI_DW 64
`define AXI_AW 32
`define AXI_NUM_MASTERS 2
`define AXI_HAS_BICMD 0
`define AXI_EN_MULTI_TILE_DLOCK_AVOID 0
`define AXI_NUM_SYS_MASTERS 2
`define AXI_NUM_SLAVES 3
`define AXI_LOG2_NS 2
`define AXI_LOG2_NM 1
`define AXI_LOG2_LCL_NMP1 2
`define AXI_LOG2_LCL_NM 1
`define AXI_LOG2_NSP1 2
`define AXI_NSP1 4
`define AXI_LOG2_NSP2 3
`define AXI_MIDW 5
`define AXI_POW2_MIDW 32
`define AXI_SIDW 6
`define AXI_BLW 8
`define AXI_HAS_TZ_SUPPORT 0
`define AXI_REMAP_EN 1
`define AXI_REMAP
`define AXI_HAS_XDCDR 0
`define AXI_TEST_XDCDR 0
`define AXI_INITIAL_LOCKDOWN 0
`define AXI_HAS_LOCKING 0
`define AXI_LOWPWR_HS_IF 0
`define AXI_LOWPWR_NOPX_CNT 32'h0
`define AXI_LOG2_LOWPWR_NOPX_CNT 1
`define AXI_INTERFACE_TYPE 1
`define AXI_HAS_AXI4 
`define AXI_HAS_QOS 0
`define AXI_DLOCK_NOTIFY_EN 0
`define AXI_DLOCK_TIMEOUT 32'd15
`define AXI_LOG2_DLOCK_TIMEOUT_P1 4
`define AXI_AR_TMO 0
`define AXI_AW_TMO 0
`define AXI_W_TMO 0
`define AXI_R_TMO 0
`define AXI_B_TMO 0
`define AXI_AR_PL_ARB 0
`define AXI_AW_PL_ARB 0
`define AXI_R_PL_ARB 0
`define AXI_W_PL_ARB 0
`define AXI_B_PL_ARB 0
`define AXI_MST_PRIORITY_W 1
`define AXI_SLV_PRIORITY_W 2
`define AXI_REG_AW_W_PATHS 1
`define AXI_MAX_UIDA 512
`define AXI_HAS_LEGAL_ADDR_OVRLP_VAL 0
`define AXI_VLD_RDY_PARITY_PROT 0
`define AXI_VLD_RDY_PARITY_MODE 0
`define AXI_HAS_EVEN_PARITY
`define IFX_RULE_SETUP 0
`define AXI_INTF_PAR_EN 0
`define AXI_INTF_PARITY_MODE 0
`define AXI_MAX_SBW 256
`define AXI_HAS_AWSB 0
`define AXI_AW_SBW 1
`define AXI_HAS_WSB 0
`define AXI_W_SBW 1
`define AXI_HAS_BSB 0
`define AXI_B_SBW 1
`define AXI_HAS_ARSB 0
`define AXI_AR_SBW 1
`define AXI_HAS_RSB 0
`define AXI_R_SBW 1
`define AXI_NV_S0_BY_M1 1
`define AXI_NV_S0_BY_M2 1
`define AXI_NV_S0_BY_M3 0
`define AXI_NV_S0_BY_M4 0
`define AXI_NV_S0_BY_M5 0
`define AXI_NV_S0_BY_M6 0
`define AXI_NV_S0_BY_M7 0
`define AXI_NV_S0_BY_M8 0
`define AXI_NV_S0_BY_M9 0
`define AXI_NV_S0_BY_M10 0
`define AXI_NV_S0_BY_M11 0
`define AXI_NV_S0_BY_M12 0
`define AXI_NV_S0_BY_M13 0
`define AXI_NV_S0_BY_M14 0
`define AXI_NV_S0_BY_M15 0
`define AXI_NV_S0_BY_M16 0
`define AXI_NV_S1_BY_M1 1
`define AXI_NV_S1_BY_M2 1
`define AXI_NV_S1_BY_M3 0
`define AXI_NV_S1_BY_M4 0
`define AXI_NV_S1_BY_M5 0
`define AXI_NV_S1_BY_M6 0
`define AXI_NV_S1_BY_M7 0
`define AXI_NV_S1_BY_M8 0
`define AXI_NV_S1_BY_M9 0
`define AXI_NV_S1_BY_M10 0
`define AXI_NV_S1_BY_M11 0
`define AXI_NV_S1_BY_M12 0
`define AXI_NV_S1_BY_M13 0
`define AXI_NV_S1_BY_M14 0
`define AXI_NV_S1_BY_M15 0
`define AXI_NV_S1_BY_M16 0
`define AXI_NV_S2_BY_M1 1
`define AXI_NV_S2_BY_M2 1
`define AXI_NV_S2_BY_M3 0
`define AXI_NV_S2_BY_M4 0
`define AXI_NV_S2_BY_M5 0
`define AXI_NV_S2_BY_M6 0
`define AXI_NV_S2_BY_M7 0
`define AXI_NV_S2_BY_M8 0
`define AXI_NV_S2_BY_M9 0
`define AXI_NV_S2_BY_M10 0
`define AXI_NV_S2_BY_M11 0
`define AXI_NV_S2_BY_M12 0
`define AXI_NV_S2_BY_M13 0
`define AXI_NV_S2_BY_M14 0
`define AXI_NV_S2_BY_M15 0
`define AXI_NV_S2_BY_M16 0
`define AXI_NV_S3_BY_M1 1
`define AXI_NV_S3_BY_M2 1
`define AXI_NV_S3_BY_M3 0
`define AXI_NV_S3_BY_M4 0
`define AXI_NV_S3_BY_M5 0
`define AXI_NV_S3_BY_M6 0
`define AXI_NV_S3_BY_M7 0
`define AXI_NV_S3_BY_M8 0
`define AXI_NV_S3_BY_M9 0
`define AXI_NV_S3_BY_M10 0
`define AXI_NV_S3_BY_M11 0
`define AXI_NV_S3_BY_M12 0
`define AXI_NV_S3_BY_M13 0
`define AXI_NV_S3_BY_M14 0
`define AXI_NV_S3_BY_M15 0
`define AXI_NV_S3_BY_M16 0
`define AXI_NV_S4_BY_M1 0
`define AXI_NV_S4_BY_M2 0
`define AXI_NV_S4_BY_M3 0
`define AXI_NV_S4_BY_M4 0
`define AXI_NV_S4_BY_M5 0
`define AXI_NV_S4_BY_M6 0
`define AXI_NV_S4_BY_M7 0
`define AXI_NV_S4_BY_M8 0
`define AXI_NV_S4_BY_M9 0
`define AXI_NV_S4_BY_M10 0
`define AXI_NV_S4_BY_M11 0
`define AXI_NV_S4_BY_M12 0
`define AXI_NV_S4_BY_M13 0
`define AXI_NV_S4_BY_M14 0
`define AXI_NV_S4_BY_M15 0
`define AXI_NV_S4_BY_M16 0
`define AXI_NV_S5_BY_M1 0
`define AXI_NV_S5_BY_M2 0
`define AXI_NV_S5_BY_M3 0
`define AXI_NV_S5_BY_M4 0
`define AXI_NV_S5_BY_M5 0
`define AXI_NV_S5_BY_M6 0
`define AXI_NV_S5_BY_M7 0
`define AXI_NV_S5_BY_M8 0
`define AXI_NV_S5_BY_M9 0
`define AXI_NV_S5_BY_M10 0
`define AXI_NV_S5_BY_M11 0
`define AXI_NV_S5_BY_M12 0
`define AXI_NV_S5_BY_M13 0
`define AXI_NV_S5_BY_M14 0
`define AXI_NV_S5_BY_M15 0
`define AXI_NV_S5_BY_M16 0
`define AXI_NV_S6_BY_M1 0
`define AXI_NV_S6_BY_M2 0
`define AXI_NV_S6_BY_M3 0
`define AXI_NV_S6_BY_M4 0
`define AXI_NV_S6_BY_M5 0
`define AXI_NV_S6_BY_M6 0
`define AXI_NV_S6_BY_M7 0
`define AXI_NV_S6_BY_M8 0
`define AXI_NV_S6_BY_M9 0
`define AXI_NV_S6_BY_M10 0
`define AXI_NV_S6_BY_M11 0
`define AXI_NV_S6_BY_M12 0
`define AXI_NV_S6_BY_M13 0
`define AXI_NV_S6_BY_M14 0
`define AXI_NV_S6_BY_M15 0
`define AXI_NV_S6_BY_M16 0
`define AXI_NV_S7_BY_M1 0
`define AXI_NV_S7_BY_M2 0
`define AXI_NV_S7_BY_M3 0
`define AXI_NV_S7_BY_M4 0
`define AXI_NV_S7_BY_M5 0
`define AXI_NV_S7_BY_M6 0
`define AXI_NV_S7_BY_M7 0
`define AXI_NV_S7_BY_M8 0
`define AXI_NV_S7_BY_M9 0
`define AXI_NV_S7_BY_M10 0
`define AXI_NV_S7_BY_M11 0
`define AXI_NV_S7_BY_M12 0
`define AXI_NV_S7_BY_M13 0
`define AXI_NV_S7_BY_M14 0
`define AXI_NV_S7_BY_M15 0
`define AXI_NV_S7_BY_M16 0
`define AXI_NV_S8_BY_M1 0
`define AXI_NV_S8_BY_M2 0
`define AXI_NV_S8_BY_M3 0
`define AXI_NV_S8_BY_M4 0
`define AXI_NV_S8_BY_M5 0
`define AXI_NV_S8_BY_M6 0
`define AXI_NV_S8_BY_M7 0
`define AXI_NV_S8_BY_M8 0
`define AXI_NV_S8_BY_M9 0
`define AXI_NV_S8_BY_M10 0
`define AXI_NV_S8_BY_M11 0
`define AXI_NV_S8_BY_M12 0
`define AXI_NV_S8_BY_M13 0
`define AXI_NV_S8_BY_M14 0
`define AXI_NV_S8_BY_M15 0
`define AXI_NV_S8_BY_M16 0
`define AXI_NV_S9_BY_M1 0
`define AXI_NV_S9_BY_M2 0
`define AXI_NV_S9_BY_M3 0
`define AXI_NV_S9_BY_M4 0
`define AXI_NV_S9_BY_M5 0
`define AXI_NV_S9_BY_M6 0
`define AXI_NV_S9_BY_M7 0
`define AXI_NV_S9_BY_M8 0
`define AXI_NV_S9_BY_M9 0
`define AXI_NV_S9_BY_M10 0
`define AXI_NV_S9_BY_M11 0
`define AXI_NV_S9_BY_M12 0
`define AXI_NV_S9_BY_M13 0
`define AXI_NV_S9_BY_M14 0
`define AXI_NV_S9_BY_M15 0
`define AXI_NV_S9_BY_M16 0
`define AXI_NV_S10_BY_M1 0
`define AXI_NV_S10_BY_M2 0
`define AXI_NV_S10_BY_M3 0
`define AXI_NV_S10_BY_M4 0
`define AXI_NV_S10_BY_M5 0
`define AXI_NV_S10_BY_M6 0
`define AXI_NV_S10_BY_M7 0
`define AXI_NV_S10_BY_M8 0
`define AXI_NV_S10_BY_M9 0
`define AXI_NV_S10_BY_M10 0
`define AXI_NV_S10_BY_M11 0
`define AXI_NV_S10_BY_M12 0
`define AXI_NV_S10_BY_M13 0
`define AXI_NV_S10_BY_M14 0
`define AXI_NV_S10_BY_M15 0
`define AXI_NV_S10_BY_M16 0
`define AXI_NV_S11_BY_M1 0
`define AXI_NV_S11_BY_M2 0
`define AXI_NV_S11_BY_M3 0
`define AXI_NV_S11_BY_M4 0
`define AXI_NV_S11_BY_M5 0
`define AXI_NV_S11_BY_M6 0
`define AXI_NV_S11_BY_M7 0
`define AXI_NV_S11_BY_M8 0
`define AXI_NV_S11_BY_M9 0
`define AXI_NV_S11_BY_M10 0
`define AXI_NV_S11_BY_M11 0
`define AXI_NV_S11_BY_M12 0
`define AXI_NV_S11_BY_M13 0
`define AXI_NV_S11_BY_M14 0
`define AXI_NV_S11_BY_M15 0
`define AXI_NV_S11_BY_M16 0
`define AXI_NV_S12_BY_M1 0
`define AXI_NV_S12_BY_M2 0
`define AXI_NV_S12_BY_M3 0
`define AXI_NV_S12_BY_M4 0
`define AXI_NV_S12_BY_M5 0
`define AXI_NV_S12_BY_M6 0
`define AXI_NV_S12_BY_M7 0
`define AXI_NV_S12_BY_M8 0
`define AXI_NV_S12_BY_M9 0
`define AXI_NV_S12_BY_M10 0
`define AXI_NV_S12_BY_M11 0
`define AXI_NV_S12_BY_M12 0
`define AXI_NV_S12_BY_M13 0
`define AXI_NV_S12_BY_M14 0
`define AXI_NV_S12_BY_M15 0
`define AXI_NV_S12_BY_M16 0
`define AXI_NV_S13_BY_M1 0
`define AXI_NV_S13_BY_M2 0
`define AXI_NV_S13_BY_M3 0
`define AXI_NV_S13_BY_M4 0
`define AXI_NV_S13_BY_M5 0
`define AXI_NV_S13_BY_M6 0
`define AXI_NV_S13_BY_M7 0
`define AXI_NV_S13_BY_M8 0
`define AXI_NV_S13_BY_M9 0
`define AXI_NV_S13_BY_M10 0
`define AXI_NV_S13_BY_M11 0
`define AXI_NV_S13_BY_M12 0
`define AXI_NV_S13_BY_M13 0
`define AXI_NV_S13_BY_M14 0
`define AXI_NV_S13_BY_M15 0
`define AXI_NV_S13_BY_M16 0
`define AXI_NV_S14_BY_M1 0
`define AXI_NV_S14_BY_M2 0
`define AXI_NV_S14_BY_M3 0
`define AXI_NV_S14_BY_M4 0
`define AXI_NV_S14_BY_M5 0
`define AXI_NV_S14_BY_M6 0
`define AXI_NV_S14_BY_M7 0
`define AXI_NV_S14_BY_M8 0
`define AXI_NV_S14_BY_M9 0
`define AXI_NV_S14_BY_M10 0
`define AXI_NV_S14_BY_M11 0
`define AXI_NV_S14_BY_M12 0
`define AXI_NV_S14_BY_M13 0
`define AXI_NV_S14_BY_M14 0
`define AXI_NV_S14_BY_M15 0
`define AXI_NV_S14_BY_M16 0
`define AXI_NV_S15_BY_M1 0
`define AXI_NV_S15_BY_M2 0
`define AXI_NV_S15_BY_M3 0
`define AXI_NV_S15_BY_M4 0
`define AXI_NV_S15_BY_M5 0
`define AXI_NV_S15_BY_M6 0
`define AXI_NV_S15_BY_M7 0
`define AXI_NV_S15_BY_M8 0
`define AXI_NV_S15_BY_M9 0
`define AXI_NV_S15_BY_M10 0
`define AXI_NV_S15_BY_M11 0
`define AXI_NV_S15_BY_M12 0
`define AXI_NV_S15_BY_M13 0
`define AXI_NV_S15_BY_M14 0
`define AXI_NV_S15_BY_M15 0
`define AXI_NV_S15_BY_M16 0
`define AXI_NV_S16_BY_M1 0
`define AXI_NV_S16_BY_M2 0
`define AXI_NV_S16_BY_M3 0
`define AXI_NV_S16_BY_M4 0
`define AXI_NV_S16_BY_M5 0
`define AXI_NV_S16_BY_M6 0
`define AXI_NV_S16_BY_M7 0
`define AXI_NV_S16_BY_M8 0
`define AXI_NV_S16_BY_M9 0
`define AXI_NV_S16_BY_M10 0
`define AXI_NV_S16_BY_M11 0
`define AXI_NV_S16_BY_M12 0
`define AXI_NV_S16_BY_M13 0
`define AXI_NV_S16_BY_M14 0
`define AXI_NV_S16_BY_M15 0
`define AXI_NV_S16_BY_M16 0
`define AXI_NV_S1_BY_ANY_M 1
`define AXI_NV_S2_BY_ANY_M 1
`define AXI_NV_S3_BY_ANY_M 1
`define AXI_NV_S4_BY_ANY_M 0
`define AXI_NV_S5_BY_ANY_M 0
`define AXI_NV_S6_BY_ANY_M 0
`define AXI_NV_S7_BY_ANY_M 0
`define AXI_NV_S8_BY_ANY_M 0
`define AXI_NV_S9_BY_ANY_M 0
`define AXI_NV_S10_BY_ANY_M 0
`define AXI_NV_S11_BY_ANY_M 0
`define AXI_NV_S12_BY_ANY_M 0
`define AXI_NV_S13_BY_ANY_M 0
`define AXI_NV_S14_BY_ANY_M 0
`define AXI_NV_S15_BY_ANY_M 0
`define AXI_NV_S16_BY_ANY_M 0
`define AXI_BV_S0_BY_M1 1
`define AXI_BV_S0_BY_M2 1
`define AXI_BV_S0_BY_M3 0
`define AXI_BV_S0_BY_M4 0
`define AXI_BV_S0_BY_M5 0
`define AXI_BV_S0_BY_M6 0
`define AXI_BV_S0_BY_M7 0
`define AXI_BV_S0_BY_M8 0
`define AXI_BV_S0_BY_M9 0
`define AXI_BV_S0_BY_M10 0
`define AXI_BV_S0_BY_M11 0
`define AXI_BV_S0_BY_M12 0
`define AXI_BV_S0_BY_M13 0
`define AXI_BV_S0_BY_M14 0
`define AXI_BV_S0_BY_M15 0
`define AXI_BV_S0_BY_M16 0
`define AXI_BV_S1_BY_M1 1
`define AXI_BV_S1_BY_M2 1
`define AXI_BV_S1_BY_M3 0
`define AXI_BV_S1_BY_M4 0
`define AXI_BV_S1_BY_M5 0
`define AXI_BV_S1_BY_M6 0
`define AXI_BV_S1_BY_M7 0
`define AXI_BV_S1_BY_M8 0
`define AXI_BV_S1_BY_M9 0
`define AXI_BV_S1_BY_M10 0
`define AXI_BV_S1_BY_M11 0
`define AXI_BV_S1_BY_M12 0
`define AXI_BV_S1_BY_M13 0
`define AXI_BV_S1_BY_M14 0
`define AXI_BV_S1_BY_M15 0
`define AXI_BV_S1_BY_M16 0
`define AXI_BV_S2_BY_M1 1
`define AXI_BV_S2_BY_M2 1
`define AXI_BV_S2_BY_M3 0
`define AXI_BV_S2_BY_M4 0
`define AXI_BV_S2_BY_M5 0
`define AXI_BV_S2_BY_M6 0
`define AXI_BV_S2_BY_M7 0
`define AXI_BV_S2_BY_M8 0
`define AXI_BV_S2_BY_M9 0
`define AXI_BV_S2_BY_M10 0
`define AXI_BV_S2_BY_M11 0
`define AXI_BV_S2_BY_M12 0
`define AXI_BV_S2_BY_M13 0
`define AXI_BV_S2_BY_M14 0
`define AXI_BV_S2_BY_M15 0
`define AXI_BV_S2_BY_M16 0
`define AXI_BV_S3_BY_M1 1
`define AXI_BV_S3_BY_M2 1
`define AXI_BV_S3_BY_M3 0
`define AXI_BV_S3_BY_M4 0
`define AXI_BV_S3_BY_M5 0
`define AXI_BV_S3_BY_M6 0
`define AXI_BV_S3_BY_M7 0
`define AXI_BV_S3_BY_M8 0
`define AXI_BV_S3_BY_M9 0
`define AXI_BV_S3_BY_M10 0
`define AXI_BV_S3_BY_M11 0
`define AXI_BV_S3_BY_M12 0
`define AXI_BV_S3_BY_M13 0
`define AXI_BV_S3_BY_M14 0
`define AXI_BV_S3_BY_M15 0
`define AXI_BV_S3_BY_M16 0
`define AXI_BV_S4_BY_M1 0
`define AXI_BV_S4_BY_M2 0
`define AXI_BV_S4_BY_M3 0
`define AXI_BV_S4_BY_M4 0
`define AXI_BV_S4_BY_M5 0
`define AXI_BV_S4_BY_M6 0
`define AXI_BV_S4_BY_M7 0
`define AXI_BV_S4_BY_M8 0
`define AXI_BV_S4_BY_M9 0
`define AXI_BV_S4_BY_M10 0
`define AXI_BV_S4_BY_M11 0
`define AXI_BV_S4_BY_M12 0
`define AXI_BV_S4_BY_M13 0
`define AXI_BV_S4_BY_M14 0
`define AXI_BV_S4_BY_M15 0
`define AXI_BV_S4_BY_M16 0
`define AXI_BV_S5_BY_M1 0
`define AXI_BV_S5_BY_M2 0
`define AXI_BV_S5_BY_M3 0
`define AXI_BV_S5_BY_M4 0
`define AXI_BV_S5_BY_M5 0
`define AXI_BV_S5_BY_M6 0
`define AXI_BV_S5_BY_M7 0
`define AXI_BV_S5_BY_M8 0
`define AXI_BV_S5_BY_M9 0
`define AXI_BV_S5_BY_M10 0
`define AXI_BV_S5_BY_M11 0
`define AXI_BV_S5_BY_M12 0
`define AXI_BV_S5_BY_M13 0
`define AXI_BV_S5_BY_M14 0
`define AXI_BV_S5_BY_M15 0
`define AXI_BV_S5_BY_M16 0
`define AXI_BV_S6_BY_M1 0
`define AXI_BV_S6_BY_M2 0
`define AXI_BV_S6_BY_M3 0
`define AXI_BV_S6_BY_M4 0
`define AXI_BV_S6_BY_M5 0
`define AXI_BV_S6_BY_M6 0
`define AXI_BV_S6_BY_M7 0
`define AXI_BV_S6_BY_M8 0
`define AXI_BV_S6_BY_M9 0
`define AXI_BV_S6_BY_M10 0
`define AXI_BV_S6_BY_M11 0
`define AXI_BV_S6_BY_M12 0
`define AXI_BV_S6_BY_M13 0
`define AXI_BV_S6_BY_M14 0
`define AXI_BV_S6_BY_M15 0
`define AXI_BV_S6_BY_M16 0
`define AXI_BV_S7_BY_M1 0
`define AXI_BV_S7_BY_M2 0
`define AXI_BV_S7_BY_M3 0
`define AXI_BV_S7_BY_M4 0
`define AXI_BV_S7_BY_M5 0
`define AXI_BV_S7_BY_M6 0
`define AXI_BV_S7_BY_M7 0
`define AXI_BV_S7_BY_M8 0
`define AXI_BV_S7_BY_M9 0
`define AXI_BV_S7_BY_M10 0
`define AXI_BV_S7_BY_M11 0
`define AXI_BV_S7_BY_M12 0
`define AXI_BV_S7_BY_M13 0
`define AXI_BV_S7_BY_M14 0
`define AXI_BV_S7_BY_M15 0
`define AXI_BV_S7_BY_M16 0
`define AXI_BV_S8_BY_M1 0
`define AXI_BV_S8_BY_M2 0
`define AXI_BV_S8_BY_M3 0
`define AXI_BV_S8_BY_M4 0
`define AXI_BV_S8_BY_M5 0
`define AXI_BV_S8_BY_M6 0
`define AXI_BV_S8_BY_M7 0
`define AXI_BV_S8_BY_M8 0
`define AXI_BV_S8_BY_M9 0
`define AXI_BV_S8_BY_M10 0
`define AXI_BV_S8_BY_M11 0
`define AXI_BV_S8_BY_M12 0
`define AXI_BV_S8_BY_M13 0
`define AXI_BV_S8_BY_M14 0
`define AXI_BV_S8_BY_M15 0
`define AXI_BV_S8_BY_M16 0
`define AXI_BV_S9_BY_M1 0
`define AXI_BV_S9_BY_M2 0
`define AXI_BV_S9_BY_M3 0
`define AXI_BV_S9_BY_M4 0
`define AXI_BV_S9_BY_M5 0
`define AXI_BV_S9_BY_M6 0
`define AXI_BV_S9_BY_M7 0
`define AXI_BV_S9_BY_M8 0
`define AXI_BV_S9_BY_M9 0
`define AXI_BV_S9_BY_M10 0
`define AXI_BV_S9_BY_M11 0
`define AXI_BV_S9_BY_M12 0
`define AXI_BV_S9_BY_M13 0
`define AXI_BV_S9_BY_M14 0
`define AXI_BV_S9_BY_M15 0
`define AXI_BV_S9_BY_M16 0
`define AXI_BV_S10_BY_M1 0
`define AXI_BV_S10_BY_M2 0
`define AXI_BV_S10_BY_M3 0
`define AXI_BV_S10_BY_M4 0
`define AXI_BV_S10_BY_M5 0
`define AXI_BV_S10_BY_M6 0
`define AXI_BV_S10_BY_M7 0
`define AXI_BV_S10_BY_M8 0
`define AXI_BV_S10_BY_M9 0
`define AXI_BV_S10_BY_M10 0
`define AXI_BV_S10_BY_M11 0
`define AXI_BV_S10_BY_M12 0
`define AXI_BV_S10_BY_M13 0
`define AXI_BV_S10_BY_M14 0
`define AXI_BV_S10_BY_M15 0
`define AXI_BV_S10_BY_M16 0
`define AXI_BV_S11_BY_M1 0
`define AXI_BV_S11_BY_M2 0
`define AXI_BV_S11_BY_M3 0
`define AXI_BV_S11_BY_M4 0
`define AXI_BV_S11_BY_M5 0
`define AXI_BV_S11_BY_M6 0
`define AXI_BV_S11_BY_M7 0
`define AXI_BV_S11_BY_M8 0
`define AXI_BV_S11_BY_M9 0
`define AXI_BV_S11_BY_M10 0
`define AXI_BV_S11_BY_M11 0
`define AXI_BV_S11_BY_M12 0
`define AXI_BV_S11_BY_M13 0
`define AXI_BV_S11_BY_M14 0
`define AXI_BV_S11_BY_M15 0
`define AXI_BV_S11_BY_M16 0
`define AXI_BV_S12_BY_M1 0
`define AXI_BV_S12_BY_M2 0
`define AXI_BV_S12_BY_M3 0
`define AXI_BV_S12_BY_M4 0
`define AXI_BV_S12_BY_M5 0
`define AXI_BV_S12_BY_M6 0
`define AXI_BV_S12_BY_M7 0
`define AXI_BV_S12_BY_M8 0
`define AXI_BV_S12_BY_M9 0
`define AXI_BV_S12_BY_M10 0
`define AXI_BV_S12_BY_M11 0
`define AXI_BV_S12_BY_M12 0
`define AXI_BV_S12_BY_M13 0
`define AXI_BV_S12_BY_M14 0
`define AXI_BV_S12_BY_M15 0
`define AXI_BV_S12_BY_M16 0
`define AXI_BV_S13_BY_M1 0
`define AXI_BV_S13_BY_M2 0
`define AXI_BV_S13_BY_M3 0
`define AXI_BV_S13_BY_M4 0
`define AXI_BV_S13_BY_M5 0
`define AXI_BV_S13_BY_M6 0
`define AXI_BV_S13_BY_M7 0
`define AXI_BV_S13_BY_M8 0
`define AXI_BV_S13_BY_M9 0
`define AXI_BV_S13_BY_M10 0
`define AXI_BV_S13_BY_M11 0
`define AXI_BV_S13_BY_M12 0
`define AXI_BV_S13_BY_M13 0
`define AXI_BV_S13_BY_M14 0
`define AXI_BV_S13_BY_M15 0
`define AXI_BV_S13_BY_M16 0
`define AXI_BV_S14_BY_M1 0
`define AXI_BV_S14_BY_M2 0
`define AXI_BV_S14_BY_M3 0
`define AXI_BV_S14_BY_M4 0
`define AXI_BV_S14_BY_M5 0
`define AXI_BV_S14_BY_M6 0
`define AXI_BV_S14_BY_M7 0
`define AXI_BV_S14_BY_M8 0
`define AXI_BV_S14_BY_M9 0
`define AXI_BV_S14_BY_M10 0
`define AXI_BV_S14_BY_M11 0
`define AXI_BV_S14_BY_M12 0
`define AXI_BV_S14_BY_M13 0
`define AXI_BV_S14_BY_M14 0
`define AXI_BV_S14_BY_M15 0
`define AXI_BV_S14_BY_M16 0
`define AXI_BV_S15_BY_M1 0
`define AXI_BV_S15_BY_M2 0
`define AXI_BV_S15_BY_M3 0
`define AXI_BV_S15_BY_M4 0
`define AXI_BV_S15_BY_M5 0
`define AXI_BV_S15_BY_M6 0
`define AXI_BV_S15_BY_M7 0
`define AXI_BV_S15_BY_M8 0
`define AXI_BV_S15_BY_M9 0
`define AXI_BV_S15_BY_M10 0
`define AXI_BV_S15_BY_M11 0
`define AXI_BV_S15_BY_M12 0
`define AXI_BV_S15_BY_M13 0
`define AXI_BV_S15_BY_M14 0
`define AXI_BV_S15_BY_M15 0
`define AXI_BV_S15_BY_M16 0
`define AXI_BV_S16_BY_M1 0
`define AXI_BV_S16_BY_M2 0
`define AXI_BV_S16_BY_M3 0
`define AXI_BV_S16_BY_M4 0
`define AXI_BV_S16_BY_M5 0
`define AXI_BV_S16_BY_M6 0
`define AXI_BV_S16_BY_M7 0
`define AXI_BV_S16_BY_M8 0
`define AXI_BV_S16_BY_M9 0
`define AXI_BV_S16_BY_M10 0
`define AXI_BV_S16_BY_M11 0
`define AXI_BV_S16_BY_M12 0
`define AXI_BV_S16_BY_M13 0
`define AXI_BV_S16_BY_M14 0
`define AXI_BV_S16_BY_M15 0
`define AXI_BV_S16_BY_M16 0
`define AXI_BV_S1_BY_ANY_M 1
`define AXI_BV_S2_BY_ANY_M 1
`define AXI_BV_S3_BY_ANY_M 1
`define AXI_BV_S4_BY_ANY_M 0
`define AXI_BV_S5_BY_ANY_M 0
`define AXI_BV_S6_BY_ANY_M 0
`define AXI_BV_S7_BY_ANY_M 0
`define AXI_BV_S8_BY_ANY_M 0
`define AXI_BV_S9_BY_ANY_M 0
`define AXI_BV_S10_BY_ANY_M 0
`define AXI_BV_S11_BY_ANY_M 0
`define AXI_BV_S12_BY_ANY_M 0
`define AXI_BV_S13_BY_ANY_M 0
`define AXI_BV_S14_BY_ANY_M 0
`define AXI_BV_S15_BY_ANY_M 0
`define AXI_BV_S16_BY_ANY_M 0
`define AXI_VV_S0_BY_M1 1
`define AXI_V_S0_BY_M1
`define AXI_VV_S0_BY_M2 1
`define AXI_V_S0_BY_M2
`define AXI_VV_S0_BY_M3 0
`define AXI_VV_S0_BY_M4 0
`define AXI_VV_S0_BY_M5 0
`define AXI_VV_S0_BY_M6 0
`define AXI_VV_S0_BY_M7 0
`define AXI_VV_S0_BY_M8 0
`define AXI_VV_S0_BY_M9 0
`define AXI_VV_S0_BY_M10 0
`define AXI_VV_S0_BY_M11 0
`define AXI_VV_S0_BY_M12 0
`define AXI_VV_S0_BY_M13 0
`define AXI_VV_S0_BY_M14 0
`define AXI_VV_S0_BY_M15 0
`define AXI_VV_S0_BY_M16 0
`define AXI_VV_S1_BY_M1 1
`define AXI_V_S1_BY_M1
`define AXI_VV_S1_BY_M2 1
`define AXI_V_S1_BY_M2
`define AXI_VV_S1_BY_M3 0
`define AXI_VV_S1_BY_M4 0
`define AXI_VV_S1_BY_M5 0
`define AXI_VV_S1_BY_M6 0
`define AXI_VV_S1_BY_M7 0
`define AXI_VV_S1_BY_M8 0
`define AXI_VV_S1_BY_M9 0
`define AXI_VV_S1_BY_M10 0
`define AXI_VV_S1_BY_M11 0
`define AXI_VV_S1_BY_M12 0
`define AXI_VV_S1_BY_M13 0
`define AXI_VV_S1_BY_M14 0
`define AXI_VV_S1_BY_M15 0
`define AXI_VV_S1_BY_M16 0
`define AXI_VV_S2_BY_M1 1
`define AXI_V_S2_BY_M1
`define AXI_VV_S2_BY_M2 1
`define AXI_V_S2_BY_M2
`define AXI_VV_S2_BY_M3 0
`define AXI_VV_S2_BY_M4 0
`define AXI_VV_S2_BY_M5 0
`define AXI_VV_S2_BY_M6 0
`define AXI_VV_S2_BY_M7 0
`define AXI_VV_S2_BY_M8 0
`define AXI_VV_S2_BY_M9 0
`define AXI_VV_S2_BY_M10 0
`define AXI_VV_S2_BY_M11 0
`define AXI_VV_S2_BY_M12 0
`define AXI_VV_S2_BY_M13 0
`define AXI_VV_S2_BY_M14 0
`define AXI_VV_S2_BY_M15 0
`define AXI_VV_S2_BY_M16 0
`define AXI_VV_S3_BY_M1 1
`define AXI_V_S3_BY_M1
`define AXI_VV_S3_BY_M2 1
`define AXI_V_S3_BY_M2
`define AXI_VV_S3_BY_M3 0
`define AXI_VV_S3_BY_M4 0
`define AXI_VV_S3_BY_M5 0
`define AXI_VV_S3_BY_M6 0
`define AXI_VV_S3_BY_M7 0
`define AXI_VV_S3_BY_M8 0
`define AXI_VV_S3_BY_M9 0
`define AXI_VV_S3_BY_M10 0
`define AXI_VV_S3_BY_M11 0
`define AXI_VV_S3_BY_M12 0
`define AXI_VV_S3_BY_M13 0
`define AXI_VV_S3_BY_M14 0
`define AXI_VV_S3_BY_M15 0
`define AXI_VV_S3_BY_M16 0
`define AXI_VV_S4_BY_M1 0
`define AXI_VV_S4_BY_M2 0
`define AXI_VV_S4_BY_M3 0
`define AXI_VV_S4_BY_M4 0
`define AXI_VV_S4_BY_M5 0
`define AXI_VV_S4_BY_M6 0
`define AXI_VV_S4_BY_M7 0
`define AXI_VV_S4_BY_M8 0
`define AXI_VV_S4_BY_M9 0
`define AXI_VV_S4_BY_M10 0
`define AXI_VV_S4_BY_M11 0
`define AXI_VV_S4_BY_M12 0
`define AXI_VV_S4_BY_M13 0
`define AXI_VV_S4_BY_M14 0
`define AXI_VV_S4_BY_M15 0
`define AXI_VV_S4_BY_M16 0
`define AXI_VV_S5_BY_M1 0
`define AXI_VV_S5_BY_M2 0
`define AXI_VV_S5_BY_M3 0
`define AXI_VV_S5_BY_M4 0
`define AXI_VV_S5_BY_M5 0
`define AXI_VV_S5_BY_M6 0
`define AXI_VV_S5_BY_M7 0
`define AXI_VV_S5_BY_M8 0
`define AXI_VV_S5_BY_M9 0
`define AXI_VV_S5_BY_M10 0
`define AXI_VV_S5_BY_M11 0
`define AXI_VV_S5_BY_M12 0
`define AXI_VV_S5_BY_M13 0
`define AXI_VV_S5_BY_M14 0
`define AXI_VV_S5_BY_M15 0
`define AXI_VV_S5_BY_M16 0
`define AXI_VV_S6_BY_M1 0
`define AXI_VV_S6_BY_M2 0
`define AXI_VV_S6_BY_M3 0
`define AXI_VV_S6_BY_M4 0
`define AXI_VV_S6_BY_M5 0
`define AXI_VV_S6_BY_M6 0
`define AXI_VV_S6_BY_M7 0
`define AXI_VV_S6_BY_M8 0
`define AXI_VV_S6_BY_M9 0
`define AXI_VV_S6_BY_M10 0
`define AXI_VV_S6_BY_M11 0
`define AXI_VV_S6_BY_M12 0
`define AXI_VV_S6_BY_M13 0
`define AXI_VV_S6_BY_M14 0
`define AXI_VV_S6_BY_M15 0
`define AXI_VV_S6_BY_M16 0
`define AXI_VV_S7_BY_M1 0
`define AXI_VV_S7_BY_M2 0
`define AXI_VV_S7_BY_M3 0
`define AXI_VV_S7_BY_M4 0
`define AXI_VV_S7_BY_M5 0
`define AXI_VV_S7_BY_M6 0
`define AXI_VV_S7_BY_M7 0
`define AXI_VV_S7_BY_M8 0
`define AXI_VV_S7_BY_M9 0
`define AXI_VV_S7_BY_M10 0
`define AXI_VV_S7_BY_M11 0
`define AXI_VV_S7_BY_M12 0
`define AXI_VV_S7_BY_M13 0
`define AXI_VV_S7_BY_M14 0
`define AXI_VV_S7_BY_M15 0
`define AXI_VV_S7_BY_M16 0
`define AXI_VV_S8_BY_M1 0
`define AXI_VV_S8_BY_M2 0
`define AXI_VV_S8_BY_M3 0
`define AXI_VV_S8_BY_M4 0
`define AXI_VV_S8_BY_M5 0
`define AXI_VV_S8_BY_M6 0
`define AXI_VV_S8_BY_M7 0
`define AXI_VV_S8_BY_M8 0
`define AXI_VV_S8_BY_M9 0
`define AXI_VV_S8_BY_M10 0
`define AXI_VV_S8_BY_M11 0
`define AXI_VV_S8_BY_M12 0
`define AXI_VV_S8_BY_M13 0
`define AXI_VV_S8_BY_M14 0
`define AXI_VV_S8_BY_M15 0
`define AXI_VV_S8_BY_M16 0
`define AXI_VV_S9_BY_M1 0
`define AXI_VV_S9_BY_M2 0
`define AXI_VV_S9_BY_M3 0
`define AXI_VV_S9_BY_M4 0
`define AXI_VV_S9_BY_M5 0
`define AXI_VV_S9_BY_M6 0
`define AXI_VV_S9_BY_M7 0
`define AXI_VV_S9_BY_M8 0
`define AXI_VV_S9_BY_M9 0
`define AXI_VV_S9_BY_M10 0
`define AXI_VV_S9_BY_M11 0
`define AXI_VV_S9_BY_M12 0
`define AXI_VV_S9_BY_M13 0
`define AXI_VV_S9_BY_M14 0
`define AXI_VV_S9_BY_M15 0
`define AXI_VV_S9_BY_M16 0
`define AXI_VV_S10_BY_M1 0
`define AXI_VV_S10_BY_M2 0
`define AXI_VV_S10_BY_M3 0
`define AXI_VV_S10_BY_M4 0
`define AXI_VV_S10_BY_M5 0
`define AXI_VV_S10_BY_M6 0
`define AXI_VV_S10_BY_M7 0
`define AXI_VV_S10_BY_M8 0
`define AXI_VV_S10_BY_M9 0
`define AXI_VV_S10_BY_M10 0
`define AXI_VV_S10_BY_M11 0
`define AXI_VV_S10_BY_M12 0
`define AXI_VV_S10_BY_M13 0
`define AXI_VV_S10_BY_M14 0
`define AXI_VV_S10_BY_M15 0
`define AXI_VV_S10_BY_M16 0
`define AXI_VV_S11_BY_M1 0
`define AXI_VV_S11_BY_M2 0
`define AXI_VV_S11_BY_M3 0
`define AXI_VV_S11_BY_M4 0
`define AXI_VV_S11_BY_M5 0
`define AXI_VV_S11_BY_M6 0
`define AXI_VV_S11_BY_M7 0
`define AXI_VV_S11_BY_M8 0
`define AXI_VV_S11_BY_M9 0
`define AXI_VV_S11_BY_M10 0
`define AXI_VV_S11_BY_M11 0
`define AXI_VV_S11_BY_M12 0
`define AXI_VV_S11_BY_M13 0
`define AXI_VV_S11_BY_M14 0
`define AXI_VV_S11_BY_M15 0
`define AXI_VV_S11_BY_M16 0
`define AXI_VV_S12_BY_M1 0
`define AXI_VV_S12_BY_M2 0
`define AXI_VV_S12_BY_M3 0
`define AXI_VV_S12_BY_M4 0
`define AXI_VV_S12_BY_M5 0
`define AXI_VV_S12_BY_M6 0
`define AXI_VV_S12_BY_M7 0
`define AXI_VV_S12_BY_M8 0
`define AXI_VV_S12_BY_M9 0
`define AXI_VV_S12_BY_M10 0
`define AXI_VV_S12_BY_M11 0
`define AXI_VV_S12_BY_M12 0
`define AXI_VV_S12_BY_M13 0
`define AXI_VV_S12_BY_M14 0
`define AXI_VV_S12_BY_M15 0
`define AXI_VV_S12_BY_M16 0
`define AXI_VV_S13_BY_M1 0
`define AXI_VV_S13_BY_M2 0
`define AXI_VV_S13_BY_M3 0
`define AXI_VV_S13_BY_M4 0
`define AXI_VV_S13_BY_M5 0
`define AXI_VV_S13_BY_M6 0
`define AXI_VV_S13_BY_M7 0
`define AXI_VV_S13_BY_M8 0
`define AXI_VV_S13_BY_M9 0
`define AXI_VV_S13_BY_M10 0
`define AXI_VV_S13_BY_M11 0
`define AXI_VV_S13_BY_M12 0
`define AXI_VV_S13_BY_M13 0
`define AXI_VV_S13_BY_M14 0
`define AXI_VV_S13_BY_M15 0
`define AXI_VV_S13_BY_M16 0
`define AXI_VV_S14_BY_M1 0
`define AXI_VV_S14_BY_M2 0
`define AXI_VV_S14_BY_M3 0
`define AXI_VV_S14_BY_M4 0
`define AXI_VV_S14_BY_M5 0
`define AXI_VV_S14_BY_M6 0
`define AXI_VV_S14_BY_M7 0
`define AXI_VV_S14_BY_M8 0
`define AXI_VV_S14_BY_M9 0
`define AXI_VV_S14_BY_M10 0
`define AXI_VV_S14_BY_M11 0
`define AXI_VV_S14_BY_M12 0
`define AXI_VV_S14_BY_M13 0
`define AXI_VV_S14_BY_M14 0
`define AXI_VV_S14_BY_M15 0
`define AXI_VV_S14_BY_M16 0
`define AXI_VV_S15_BY_M1 0
`define AXI_VV_S15_BY_M2 0
`define AXI_VV_S15_BY_M3 0
`define AXI_VV_S15_BY_M4 0
`define AXI_VV_S15_BY_M5 0
`define AXI_VV_S15_BY_M6 0
`define AXI_VV_S15_BY_M7 0
`define AXI_VV_S15_BY_M8 0
`define AXI_VV_S15_BY_M9 0
`define AXI_VV_S15_BY_M10 0
`define AXI_VV_S15_BY_M11 0
`define AXI_VV_S15_BY_M12 0
`define AXI_VV_S15_BY_M13 0
`define AXI_VV_S15_BY_M14 0
`define AXI_VV_S15_BY_M15 0
`define AXI_VV_S15_BY_M16 0
`define AXI_VV_S16_BY_M1 0
`define AXI_VV_S16_BY_M2 0
`define AXI_VV_S16_BY_M3 0
`define AXI_VV_S16_BY_M4 0
`define AXI_VV_S16_BY_M5 0
`define AXI_VV_S16_BY_M6 0
`define AXI_VV_S16_BY_M7 0
`define AXI_VV_S16_BY_M8 0
`define AXI_VV_S16_BY_M9 0
`define AXI_VV_S16_BY_M10 0
`define AXI_VV_S16_BY_M11 0
`define AXI_VV_S16_BY_M12 0
`define AXI_VV_S16_BY_M13 0
`define AXI_VV_S16_BY_M14 0
`define AXI_VV_S16_BY_M15 0
`define AXI_VV_S16_BY_M16 0
`define AXI_NMV_S1 2
`define AXI_LOG2_NMV_S1 1
`define AXI_LOG2_NMP1V_S1 2
`define AXI_NMV_S2 2
`define AXI_LOG2_NMV_S2 1
`define AXI_LOG2_NMP1V_S2 2
`define AXI_NMV_S3 2
`define AXI_LOG2_NMV_S3 1
`define AXI_LOG2_NMP1V_S3 2
`define AXI_NMV_S4 1
`define AXI_LOG2_NMV_S4 1
`define AXI_LOG2_NMP1V_S4 1
`define AXI_NMV_S5 1
`define AXI_LOG2_NMV_S5 1
`define AXI_LOG2_NMP1V_S5 1
`define AXI_NMV_S6 1
`define AXI_LOG2_NMV_S6 1
`define AXI_LOG2_NMP1V_S6 1
`define AXI_NMV_S7 1
`define AXI_LOG2_NMV_S7 1
`define AXI_LOG2_NMP1V_S7 1
`define AXI_NMV_S8 1
`define AXI_LOG2_NMV_S8 1
`define AXI_LOG2_NMP1V_S8 1
`define AXI_NMV_S9 1
`define AXI_LOG2_NMV_S9 1
`define AXI_LOG2_NMP1V_S9 1
`define AXI_NMV_S10 1
`define AXI_LOG2_NMV_S10 1
`define AXI_LOG2_NMP1V_S10 1
`define AXI_NMV_S11 1
`define AXI_LOG2_NMV_S11 1
`define AXI_LOG2_NMP1V_S11 1
`define AXI_NMV_S12 1
`define AXI_LOG2_NMV_S12 1
`define AXI_LOG2_NMP1V_S12 1
`define AXI_NMV_S13 1
`define AXI_LOG2_NMV_S13 1
`define AXI_LOG2_NMP1V_S13 1
`define AXI_NMV_S14 1
`define AXI_LOG2_NMV_S14 1
`define AXI_LOG2_NMP1V_S14 1
`define AXI_NMV_S15 1
`define AXI_LOG2_NMV_S15 1
`define AXI_LOG2_NMP1V_S15 1
`define AXI_NMV_S16 1
`define AXI_LOG2_NMV_S16 1
`define AXI_LOG2_NMP1V_S16 1
`define AXI_NSV_M1 3
`define AXI_LOG2_NSV_M1 2
`define AXI_NSV_M2 3
`define AXI_LOG2_NSV_M2 2
`define AXI_NSV_M3 1
`define AXI_LOG2_NSV_M3 1
`define AXI_NSV_M4 1
`define AXI_LOG2_NSV_M4 1
`define AXI_NSV_M5 1
`define AXI_LOG2_NSV_M5 1
`define AXI_NSV_M6 1
`define AXI_LOG2_NSV_M6 1
`define AXI_NSV_M7 1
`define AXI_LOG2_NSV_M7 1
`define AXI_NSV_M8 1
`define AXI_LOG2_NSV_M8 1
`define AXI_NSV_M9 1
`define AXI_LOG2_NSV_M9 1
`define AXI_NSV_M10 1
`define AXI_LOG2_NSV_M10 1
`define AXI_NSV_M11 1
`define AXI_LOG2_NSV_M11 1
`define AXI_NSV_M12 1
`define AXI_LOG2_NSV_M12 1
`define AXI_NSV_M13 1
`define AXI_LOG2_NSV_M13 1
`define AXI_NSV_M14 1
`define AXI_LOG2_NSV_M14 1
`define AXI_NSV_M15 1
`define AXI_LOG2_NSV_M15 1
`define AXI_NSV_M16 1
`define AXI_LOG2_NSV_M16 1
`define AXI_NNMV_S1 2
`define AXI_BNMV_S1 2
`define AXI_NNMV_S2 2
`define AXI_BNMV_S2 2
`define AXI_NNMV_S3 2
`define AXI_BNMV_S3 2
`define AXI_NNMV_S4 0
`define AXI_BNMV_S4 0
`define AXI_NNMV_S5 0
`define AXI_BNMV_S5 0
`define AXI_NNMV_S6 0
`define AXI_BNMV_S6 0
`define AXI_NNMV_S7 0
`define AXI_BNMV_S7 0
`define AXI_NNMV_S8 0
`define AXI_BNMV_S8 0
`define AXI_NNMV_S9 0
`define AXI_BNMV_S9 0
`define AXI_NNMV_S10 0
`define AXI_BNMV_S10 0
`define AXI_NNMV_S11 0
`define AXI_BNMV_S11 0
`define AXI_NNMV_S12 0
`define AXI_BNMV_S12 0
`define AXI_NNMV_S13 0
`define AXI_BNMV_S13 0
`define AXI_NNMV_S14 0
`define AXI_BNMV_S14 0
`define AXI_NNMV_S15 0
`define AXI_BNMV_S15 0
`define AXI_NNMV_S16 0
`define AXI_BNMV_S16 0
`define AXI_NSP1V_M1 4
`define AXI_LOG2_NSP1V_M1 2
`define AXI_LOG2_NSP2V_M1 3
`define AXI_NSP1V_M2 4
`define AXI_LOG2_NSP1V_M2 2
`define AXI_LOG2_NSP2V_M2 3
`define AXI_NSP1V_M3 1
`define AXI_LOG2_NSP1V_M3 1
`define AXI_LOG2_NSP2V_M3 2
`define AXI_NSP1V_M4 1
`define AXI_LOG2_NSP1V_M4 1
`define AXI_LOG2_NSP2V_M4 2
`define AXI_NSP1V_M5 1
`define AXI_LOG2_NSP1V_M5 1
`define AXI_LOG2_NSP2V_M5 2
`define AXI_NSP1V_M6 1
`define AXI_LOG2_NSP1V_M6 1
`define AXI_LOG2_NSP2V_M6 2
`define AXI_NSP1V_M7 1
`define AXI_LOG2_NSP1V_M7 1
`define AXI_LOG2_NSP2V_M7 2
`define AXI_NSP1V_M8 1
`define AXI_LOG2_NSP1V_M8 1
`define AXI_LOG2_NSP2V_M8 2
`define AXI_NSP1V_M9 1
`define AXI_LOG2_NSP1V_M9 1
`define AXI_LOG2_NSP2V_M9 2
`define AXI_NSP1V_M10 1
`define AXI_LOG2_NSP1V_M10 1
`define AXI_LOG2_NSP2V_M10 2
`define AXI_NSP1V_M11 1
`define AXI_LOG2_NSP1V_M11 1
`define AXI_LOG2_NSP2V_M11 2
`define AXI_NSP1V_M12 1
`define AXI_LOG2_NSP1V_M12 1
`define AXI_LOG2_NSP2V_M12 2
`define AXI_NSP1V_M13 1
`define AXI_LOG2_NSP1V_M13 1
`define AXI_LOG2_NSP2V_M13 2
`define AXI_NSP1V_M14 1
`define AXI_LOG2_NSP1V_M14 1
`define AXI_LOG2_NSP2V_M14 2
`define AXI_NSP1V_M15 1
`define AXI_LOG2_NSP1V_M15 1
`define AXI_LOG2_NSP2V_M15 2
`define AXI_NSP1V_M16 1
`define AXI_LOG2_NSP1V_M16 1
`define AXI_LOG2_NSP2V_M16 2
`define AXI_ALL_AR_LAYER_SHARED 0
`define AXI_AR_LAYER_S0_M1 0
`define AXI_AR_LAYER_S0_M2 0
`define AXI_AR_LAYER_S0_M3 0
`define AXI_AR_LAYER_S0_M4 0
`define AXI_AR_LAYER_S0_M5 0
`define AXI_AR_LAYER_S0_M6 0
`define AXI_AR_LAYER_S0_M7 0
`define AXI_AR_LAYER_S0_M8 0
`define AXI_AR_LAYER_S0_M9 0
`define AXI_AR_LAYER_S0_M10 0
`define AXI_AR_LAYER_S0_M11 0
`define AXI_AR_LAYER_S0_M12 0
`define AXI_AR_LAYER_S0_M13 0
`define AXI_AR_LAYER_S0_M14 0
`define AXI_AR_LAYER_S0_M15 0
`define AXI_AR_LAYER_S0_M16 0
`define AXI_ALL_AW_LAYER_SHARED 0
`define AXI_AW_LAYER_S0_M1 0
`define AXI_AW_LAYER_S0_M2 0
`define AXI_AW_LAYER_S0_M3 0
`define AXI_AW_LAYER_S0_M4 0
`define AXI_AW_LAYER_S0_M5 0
`define AXI_AW_LAYER_S0_M6 0
`define AXI_AW_LAYER_S0_M7 0
`define AXI_AW_LAYER_S0_M8 0
`define AXI_AW_LAYER_S0_M9 0
`define AXI_AW_LAYER_S0_M10 0
`define AXI_AW_LAYER_S0_M11 0
`define AXI_AW_LAYER_S0_M12 0
`define AXI_AW_LAYER_S0_M13 0
`define AXI_AW_LAYER_S0_M14 0
`define AXI_AW_LAYER_S0_M15 0
`define AXI_AW_LAYER_S0_M16 0
`define AXI_ALL_W_LAYER_SHARED 0
`define AXI_W_LAYER_S0_M1 0
`define AXI_W_LAYER_S0_M2 0
`define AXI_W_LAYER_S0_M3 0
`define AXI_W_LAYER_S0_M4 0
`define AXI_W_LAYER_S0_M5 0
`define AXI_W_LAYER_S0_M6 0
`define AXI_W_LAYER_S0_M7 0
`define AXI_W_LAYER_S0_M8 0
`define AXI_W_LAYER_S0_M9 0
`define AXI_W_LAYER_S0_M10 0
`define AXI_W_LAYER_S0_M11 0
`define AXI_W_LAYER_S0_M12 0
`define AXI_W_LAYER_S0_M13 0
`define AXI_W_LAYER_S0_M14 0
`define AXI_W_LAYER_S0_M15 0
`define AXI_W_LAYER_S0_M16 0
`define AXI_AR_LAYER_S1_M1 0
`define AXI_AR_LAYER_S1_M2 0
`define AXI_AR_LAYER_S1_M3 0
`define AXI_AR_LAYER_S1_M4 0
`define AXI_AR_LAYER_S1_M5 0
`define AXI_AR_LAYER_S1_M6 0
`define AXI_AR_LAYER_S1_M7 0
`define AXI_AR_LAYER_S1_M8 0
`define AXI_AR_LAYER_S1_M9 0
`define AXI_AR_LAYER_S1_M10 0
`define AXI_AR_LAYER_S1_M11 0
`define AXI_AR_LAYER_S1_M12 0
`define AXI_AR_LAYER_S1_M13 0
`define AXI_AR_LAYER_S1_M14 0
`define AXI_AR_LAYER_S1_M15 0
`define AXI_AR_LAYER_S1_M16 0
`define AXI_AW_LAYER_S1_M1 0
`define AXI_AW_LAYER_S1_M2 0
`define AXI_AW_LAYER_S1_M3 0
`define AXI_AW_LAYER_S1_M4 0
`define AXI_AW_LAYER_S1_M5 0
`define AXI_AW_LAYER_S1_M6 0
`define AXI_AW_LAYER_S1_M7 0
`define AXI_AW_LAYER_S1_M8 0
`define AXI_AW_LAYER_S1_M9 0
`define AXI_AW_LAYER_S1_M10 0
`define AXI_AW_LAYER_S1_M11 0
`define AXI_AW_LAYER_S1_M12 0
`define AXI_AW_LAYER_S1_M13 0
`define AXI_AW_LAYER_S1_M14 0
`define AXI_AW_LAYER_S1_M15 0
`define AXI_AW_LAYER_S1_M16 0
`define AXI_W_LAYER_S1_M1 0
`define AXI_W_LAYER_S1_M2 0
`define AXI_W_LAYER_S1_M3 0
`define AXI_W_LAYER_S1_M4 0
`define AXI_W_LAYER_S1_M5 0
`define AXI_W_LAYER_S1_M6 0
`define AXI_W_LAYER_S1_M7 0
`define AXI_W_LAYER_S1_M8 0
`define AXI_W_LAYER_S1_M9 0
`define AXI_W_LAYER_S1_M10 0
`define AXI_W_LAYER_S1_M11 0
`define AXI_W_LAYER_S1_M12 0
`define AXI_W_LAYER_S1_M13 0
`define AXI_W_LAYER_S1_M14 0
`define AXI_W_LAYER_S1_M15 0
`define AXI_W_LAYER_S1_M16 0
`define AXI_AR_LAYER_S2_M1 0
`define AXI_AR_LAYER_S2_M2 0
`define AXI_AR_LAYER_S2_M3 0
`define AXI_AR_LAYER_S2_M4 0
`define AXI_AR_LAYER_S2_M5 0
`define AXI_AR_LAYER_S2_M6 0
`define AXI_AR_LAYER_S2_M7 0
`define AXI_AR_LAYER_S2_M8 0
`define AXI_AR_LAYER_S2_M9 0
`define AXI_AR_LAYER_S2_M10 0
`define AXI_AR_LAYER_S2_M11 0
`define AXI_AR_LAYER_S2_M12 0
`define AXI_AR_LAYER_S2_M13 0
`define AXI_AR_LAYER_S2_M14 0
`define AXI_AR_LAYER_S2_M15 0
`define AXI_AR_LAYER_S2_M16 0
`define AXI_AW_LAYER_S2_M1 0
`define AXI_AW_LAYER_S2_M2 0
`define AXI_AW_LAYER_S2_M3 0
`define AXI_AW_LAYER_S2_M4 0
`define AXI_AW_LAYER_S2_M5 0
`define AXI_AW_LAYER_S2_M6 0
`define AXI_AW_LAYER_S2_M7 0
`define AXI_AW_LAYER_S2_M8 0
`define AXI_AW_LAYER_S2_M9 0
`define AXI_AW_LAYER_S2_M10 0
`define AXI_AW_LAYER_S2_M11 0
`define AXI_AW_LAYER_S2_M12 0
`define AXI_AW_LAYER_S2_M13 0
`define AXI_AW_LAYER_S2_M14 0
`define AXI_AW_LAYER_S2_M15 0
`define AXI_AW_LAYER_S2_M16 0
`define AXI_W_LAYER_S2_M1 0
`define AXI_W_LAYER_S2_M2 0
`define AXI_W_LAYER_S2_M3 0
`define AXI_W_LAYER_S2_M4 0
`define AXI_W_LAYER_S2_M5 0
`define AXI_W_LAYER_S2_M6 0
`define AXI_W_LAYER_S2_M7 0
`define AXI_W_LAYER_S2_M8 0
`define AXI_W_LAYER_S2_M9 0
`define AXI_W_LAYER_S2_M10 0
`define AXI_W_LAYER_S2_M11 0
`define AXI_W_LAYER_S2_M12 0
`define AXI_W_LAYER_S2_M13 0
`define AXI_W_LAYER_S2_M14 0
`define AXI_W_LAYER_S2_M15 0
`define AXI_W_LAYER_S2_M16 0
`define AXI_AR_LAYER_S3_M1 0
`define AXI_AR_LAYER_S3_M2 0
`define AXI_AR_LAYER_S3_M3 0
`define AXI_AR_LAYER_S3_M4 0
`define AXI_AR_LAYER_S3_M5 0
`define AXI_AR_LAYER_S3_M6 0
`define AXI_AR_LAYER_S3_M7 0
`define AXI_AR_LAYER_S3_M8 0
`define AXI_AR_LAYER_S3_M9 0
`define AXI_AR_LAYER_S3_M10 0
`define AXI_AR_LAYER_S3_M11 0
`define AXI_AR_LAYER_S3_M12 0
`define AXI_AR_LAYER_S3_M13 0
`define AXI_AR_LAYER_S3_M14 0
`define AXI_AR_LAYER_S3_M15 0
`define AXI_AR_LAYER_S3_M16 0
`define AXI_AW_LAYER_S3_M1 0
`define AXI_AW_LAYER_S3_M2 0
`define AXI_AW_LAYER_S3_M3 0
`define AXI_AW_LAYER_S3_M4 0
`define AXI_AW_LAYER_S3_M5 0
`define AXI_AW_LAYER_S3_M6 0
`define AXI_AW_LAYER_S3_M7 0
`define AXI_AW_LAYER_S3_M8 0
`define AXI_AW_LAYER_S3_M9 0
`define AXI_AW_LAYER_S3_M10 0
`define AXI_AW_LAYER_S3_M11 0
`define AXI_AW_LAYER_S3_M12 0
`define AXI_AW_LAYER_S3_M13 0
`define AXI_AW_LAYER_S3_M14 0
`define AXI_AW_LAYER_S3_M15 0
`define AXI_AW_LAYER_S3_M16 0
`define AXI_W_LAYER_S3_M1 0
`define AXI_W_LAYER_S3_M2 0
`define AXI_W_LAYER_S3_M3 0
`define AXI_W_LAYER_S3_M4 0
`define AXI_W_LAYER_S3_M5 0
`define AXI_W_LAYER_S3_M6 0
`define AXI_W_LAYER_S3_M7 0
`define AXI_W_LAYER_S3_M8 0
`define AXI_W_LAYER_S3_M9 0
`define AXI_W_LAYER_S3_M10 0
`define AXI_W_LAYER_S3_M11 0
`define AXI_W_LAYER_S3_M12 0
`define AXI_W_LAYER_S3_M13 0
`define AXI_W_LAYER_S3_M14 0
`define AXI_W_LAYER_S3_M15 0
`define AXI_W_LAYER_S3_M16 0
`define AXI_AR_LAYER_S4_M1 0
`define AXI_AR_LAYER_S4_M2 0
`define AXI_AR_LAYER_S4_M3 0
`define AXI_AR_LAYER_S4_M4 0
`define AXI_AR_LAYER_S4_M5 0
`define AXI_AR_LAYER_S4_M6 0
`define AXI_AR_LAYER_S4_M7 0
`define AXI_AR_LAYER_S4_M8 0
`define AXI_AR_LAYER_S4_M9 0
`define AXI_AR_LAYER_S4_M10 0
`define AXI_AR_LAYER_S4_M11 0
`define AXI_AR_LAYER_S4_M12 0
`define AXI_AR_LAYER_S4_M13 0
`define AXI_AR_LAYER_S4_M14 0
`define AXI_AR_LAYER_S4_M15 0
`define AXI_AR_LAYER_S4_M16 0
`define AXI_AW_LAYER_S4_M1 0
`define AXI_AW_LAYER_S4_M2 0
`define AXI_AW_LAYER_S4_M3 0
`define AXI_AW_LAYER_S4_M4 0
`define AXI_AW_LAYER_S4_M5 0
`define AXI_AW_LAYER_S4_M6 0
`define AXI_AW_LAYER_S4_M7 0
`define AXI_AW_LAYER_S4_M8 0
`define AXI_AW_LAYER_S4_M9 0
`define AXI_AW_LAYER_S4_M10 0
`define AXI_AW_LAYER_S4_M11 0
`define AXI_AW_LAYER_S4_M12 0
`define AXI_AW_LAYER_S4_M13 0
`define AXI_AW_LAYER_S4_M14 0
`define AXI_AW_LAYER_S4_M15 0
`define AXI_AW_LAYER_S4_M16 0
`define AXI_W_LAYER_S4_M1 0
`define AXI_W_LAYER_S4_M2 0
`define AXI_W_LAYER_S4_M3 0
`define AXI_W_LAYER_S4_M4 0
`define AXI_W_LAYER_S4_M5 0
`define AXI_W_LAYER_S4_M6 0
`define AXI_W_LAYER_S4_M7 0
`define AXI_W_LAYER_S4_M8 0
`define AXI_W_LAYER_S4_M9 0
`define AXI_W_LAYER_S4_M10 0
`define AXI_W_LAYER_S4_M11 0
`define AXI_W_LAYER_S4_M12 0
`define AXI_W_LAYER_S4_M13 0
`define AXI_W_LAYER_S4_M14 0
`define AXI_W_LAYER_S4_M15 0
`define AXI_W_LAYER_S4_M16 0
`define AXI_AR_LAYER_S5_M1 0
`define AXI_AR_LAYER_S5_M2 0
`define AXI_AR_LAYER_S5_M3 0
`define AXI_AR_LAYER_S5_M4 0
`define AXI_AR_LAYER_S5_M5 0
`define AXI_AR_LAYER_S5_M6 0
`define AXI_AR_LAYER_S5_M7 0
`define AXI_AR_LAYER_S5_M8 0
`define AXI_AR_LAYER_S5_M9 0
`define AXI_AR_LAYER_S5_M10 0
`define AXI_AR_LAYER_S5_M11 0
`define AXI_AR_LAYER_S5_M12 0
`define AXI_AR_LAYER_S5_M13 0
`define AXI_AR_LAYER_S5_M14 0
`define AXI_AR_LAYER_S5_M15 0
`define AXI_AR_LAYER_S5_M16 0
`define AXI_AW_LAYER_S5_M1 0
`define AXI_AW_LAYER_S5_M2 0
`define AXI_AW_LAYER_S5_M3 0
`define AXI_AW_LAYER_S5_M4 0
`define AXI_AW_LAYER_S5_M5 0
`define AXI_AW_LAYER_S5_M6 0
`define AXI_AW_LAYER_S5_M7 0
`define AXI_AW_LAYER_S5_M8 0
`define AXI_AW_LAYER_S5_M9 0
`define AXI_AW_LAYER_S5_M10 0
`define AXI_AW_LAYER_S5_M11 0
`define AXI_AW_LAYER_S5_M12 0
`define AXI_AW_LAYER_S5_M13 0
`define AXI_AW_LAYER_S5_M14 0
`define AXI_AW_LAYER_S5_M15 0
`define AXI_AW_LAYER_S5_M16 0
`define AXI_W_LAYER_S5_M1 0
`define AXI_W_LAYER_S5_M2 0
`define AXI_W_LAYER_S5_M3 0
`define AXI_W_LAYER_S5_M4 0
`define AXI_W_LAYER_S5_M5 0
`define AXI_W_LAYER_S5_M6 0
`define AXI_W_LAYER_S5_M7 0
`define AXI_W_LAYER_S5_M8 0
`define AXI_W_LAYER_S5_M9 0
`define AXI_W_LAYER_S5_M10 0
`define AXI_W_LAYER_S5_M11 0
`define AXI_W_LAYER_S5_M12 0
`define AXI_W_LAYER_S5_M13 0
`define AXI_W_LAYER_S5_M14 0
`define AXI_W_LAYER_S5_M15 0
`define AXI_W_LAYER_S5_M16 0
`define AXI_AR_LAYER_S6_M1 0
`define AXI_AR_LAYER_S6_M2 0
`define AXI_AR_LAYER_S6_M3 0
`define AXI_AR_LAYER_S6_M4 0
`define AXI_AR_LAYER_S6_M5 0
`define AXI_AR_LAYER_S6_M6 0
`define AXI_AR_LAYER_S6_M7 0
`define AXI_AR_LAYER_S6_M8 0
`define AXI_AR_LAYER_S6_M9 0
`define AXI_AR_LAYER_S6_M10 0
`define AXI_AR_LAYER_S6_M11 0
`define AXI_AR_LAYER_S6_M12 0
`define AXI_AR_LAYER_S6_M13 0
`define AXI_AR_LAYER_S6_M14 0
`define AXI_AR_LAYER_S6_M15 0
`define AXI_AR_LAYER_S6_M16 0
`define AXI_AW_LAYER_S6_M1 0
`define AXI_AW_LAYER_S6_M2 0
`define AXI_AW_LAYER_S6_M3 0
`define AXI_AW_LAYER_S6_M4 0
`define AXI_AW_LAYER_S6_M5 0
`define AXI_AW_LAYER_S6_M6 0
`define AXI_AW_LAYER_S6_M7 0
`define AXI_AW_LAYER_S6_M8 0
`define AXI_AW_LAYER_S6_M9 0
`define AXI_AW_LAYER_S6_M10 0
`define AXI_AW_LAYER_S6_M11 0
`define AXI_AW_LAYER_S6_M12 0
`define AXI_AW_LAYER_S6_M13 0
`define AXI_AW_LAYER_S6_M14 0
`define AXI_AW_LAYER_S6_M15 0
`define AXI_AW_LAYER_S6_M16 0
`define AXI_W_LAYER_S6_M1 0
`define AXI_W_LAYER_S6_M2 0
`define AXI_W_LAYER_S6_M3 0
`define AXI_W_LAYER_S6_M4 0
`define AXI_W_LAYER_S6_M5 0
`define AXI_W_LAYER_S6_M6 0
`define AXI_W_LAYER_S6_M7 0
`define AXI_W_LAYER_S6_M8 0
`define AXI_W_LAYER_S6_M9 0
`define AXI_W_LAYER_S6_M10 0
`define AXI_W_LAYER_S6_M11 0
`define AXI_W_LAYER_S6_M12 0
`define AXI_W_LAYER_S6_M13 0
`define AXI_W_LAYER_S6_M14 0
`define AXI_W_LAYER_S6_M15 0
`define AXI_W_LAYER_S6_M16 0
`define AXI_AR_LAYER_S7_M1 0
`define AXI_AR_LAYER_S7_M2 0
`define AXI_AR_LAYER_S7_M3 0
`define AXI_AR_LAYER_S7_M4 0
`define AXI_AR_LAYER_S7_M5 0
`define AXI_AR_LAYER_S7_M6 0
`define AXI_AR_LAYER_S7_M7 0
`define AXI_AR_LAYER_S7_M8 0
`define AXI_AR_LAYER_S7_M9 0
`define AXI_AR_LAYER_S7_M10 0
`define AXI_AR_LAYER_S7_M11 0
`define AXI_AR_LAYER_S7_M12 0
`define AXI_AR_LAYER_S7_M13 0
`define AXI_AR_LAYER_S7_M14 0
`define AXI_AR_LAYER_S7_M15 0
`define AXI_AR_LAYER_S7_M16 0
`define AXI_AW_LAYER_S7_M1 0
`define AXI_AW_LAYER_S7_M2 0
`define AXI_AW_LAYER_S7_M3 0
`define AXI_AW_LAYER_S7_M4 0
`define AXI_AW_LAYER_S7_M5 0
`define AXI_AW_LAYER_S7_M6 0
`define AXI_AW_LAYER_S7_M7 0
`define AXI_AW_LAYER_S7_M8 0
`define AXI_AW_LAYER_S7_M9 0
`define AXI_AW_LAYER_S7_M10 0
`define AXI_AW_LAYER_S7_M11 0
`define AXI_AW_LAYER_S7_M12 0
`define AXI_AW_LAYER_S7_M13 0
`define AXI_AW_LAYER_S7_M14 0
`define AXI_AW_LAYER_S7_M15 0
`define AXI_AW_LAYER_S7_M16 0
`define AXI_W_LAYER_S7_M1 0
`define AXI_W_LAYER_S7_M2 0
`define AXI_W_LAYER_S7_M3 0
`define AXI_W_LAYER_S7_M4 0
`define AXI_W_LAYER_S7_M5 0
`define AXI_W_LAYER_S7_M6 0
`define AXI_W_LAYER_S7_M7 0
`define AXI_W_LAYER_S7_M8 0
`define AXI_W_LAYER_S7_M9 0
`define AXI_W_LAYER_S7_M10 0
`define AXI_W_LAYER_S7_M11 0
`define AXI_W_LAYER_S7_M12 0
`define AXI_W_LAYER_S7_M13 0
`define AXI_W_LAYER_S7_M14 0
`define AXI_W_LAYER_S7_M15 0
`define AXI_W_LAYER_S7_M16 0
`define AXI_AR_LAYER_S8_M1 0
`define AXI_AR_LAYER_S8_M2 0
`define AXI_AR_LAYER_S8_M3 0
`define AXI_AR_LAYER_S8_M4 0
`define AXI_AR_LAYER_S8_M5 0
`define AXI_AR_LAYER_S8_M6 0
`define AXI_AR_LAYER_S8_M7 0
`define AXI_AR_LAYER_S8_M8 0
`define AXI_AR_LAYER_S8_M9 0
`define AXI_AR_LAYER_S8_M10 0
`define AXI_AR_LAYER_S8_M11 0
`define AXI_AR_LAYER_S8_M12 0
`define AXI_AR_LAYER_S8_M13 0
`define AXI_AR_LAYER_S8_M14 0
`define AXI_AR_LAYER_S8_M15 0
`define AXI_AR_LAYER_S8_M16 0
`define AXI_AW_LAYER_S8_M1 0
`define AXI_AW_LAYER_S8_M2 0
`define AXI_AW_LAYER_S8_M3 0
`define AXI_AW_LAYER_S8_M4 0
`define AXI_AW_LAYER_S8_M5 0
`define AXI_AW_LAYER_S8_M6 0
`define AXI_AW_LAYER_S8_M7 0
`define AXI_AW_LAYER_S8_M8 0
`define AXI_AW_LAYER_S8_M9 0
`define AXI_AW_LAYER_S8_M10 0
`define AXI_AW_LAYER_S8_M11 0
`define AXI_AW_LAYER_S8_M12 0
`define AXI_AW_LAYER_S8_M13 0
`define AXI_AW_LAYER_S8_M14 0
`define AXI_AW_LAYER_S8_M15 0
`define AXI_AW_LAYER_S8_M16 0
`define AXI_W_LAYER_S8_M1 0
`define AXI_W_LAYER_S8_M2 0
`define AXI_W_LAYER_S8_M3 0
`define AXI_W_LAYER_S8_M4 0
`define AXI_W_LAYER_S8_M5 0
`define AXI_W_LAYER_S8_M6 0
`define AXI_W_LAYER_S8_M7 0
`define AXI_W_LAYER_S8_M8 0
`define AXI_W_LAYER_S8_M9 0
`define AXI_W_LAYER_S8_M10 0
`define AXI_W_LAYER_S8_M11 0
`define AXI_W_LAYER_S8_M12 0
`define AXI_W_LAYER_S8_M13 0
`define AXI_W_LAYER_S8_M14 0
`define AXI_W_LAYER_S8_M15 0
`define AXI_W_LAYER_S8_M16 0
`define AXI_AR_LAYER_S9_M1 0
`define AXI_AR_LAYER_S9_M2 0
`define AXI_AR_LAYER_S9_M3 0
`define AXI_AR_LAYER_S9_M4 0
`define AXI_AR_LAYER_S9_M5 0
`define AXI_AR_LAYER_S9_M6 0
`define AXI_AR_LAYER_S9_M7 0
`define AXI_AR_LAYER_S9_M8 0
`define AXI_AR_LAYER_S9_M9 0
`define AXI_AR_LAYER_S9_M10 0
`define AXI_AR_LAYER_S9_M11 0
`define AXI_AR_LAYER_S9_M12 0
`define AXI_AR_LAYER_S9_M13 0
`define AXI_AR_LAYER_S9_M14 0
`define AXI_AR_LAYER_S9_M15 0
`define AXI_AR_LAYER_S9_M16 0
`define AXI_AW_LAYER_S9_M1 0
`define AXI_AW_LAYER_S9_M2 0
`define AXI_AW_LAYER_S9_M3 0
`define AXI_AW_LAYER_S9_M4 0
`define AXI_AW_LAYER_S9_M5 0
`define AXI_AW_LAYER_S9_M6 0
`define AXI_AW_LAYER_S9_M7 0
`define AXI_AW_LAYER_S9_M8 0
`define AXI_AW_LAYER_S9_M9 0
`define AXI_AW_LAYER_S9_M10 0
`define AXI_AW_LAYER_S9_M11 0
`define AXI_AW_LAYER_S9_M12 0
`define AXI_AW_LAYER_S9_M13 0
`define AXI_AW_LAYER_S9_M14 0
`define AXI_AW_LAYER_S9_M15 0
`define AXI_AW_LAYER_S9_M16 0
`define AXI_W_LAYER_S9_M1 0
`define AXI_W_LAYER_S9_M2 0
`define AXI_W_LAYER_S9_M3 0
`define AXI_W_LAYER_S9_M4 0
`define AXI_W_LAYER_S9_M5 0
`define AXI_W_LAYER_S9_M6 0
`define AXI_W_LAYER_S9_M7 0
`define AXI_W_LAYER_S9_M8 0
`define AXI_W_LAYER_S9_M9 0
`define AXI_W_LAYER_S9_M10 0
`define AXI_W_LAYER_S9_M11 0
`define AXI_W_LAYER_S9_M12 0
`define AXI_W_LAYER_S9_M13 0
`define AXI_W_LAYER_S9_M14 0
`define AXI_W_LAYER_S9_M15 0
`define AXI_W_LAYER_S9_M16 0
`define AXI_AR_LAYER_S10_M1 0
`define AXI_AR_LAYER_S10_M2 0
`define AXI_AR_LAYER_S10_M3 0
`define AXI_AR_LAYER_S10_M4 0
`define AXI_AR_LAYER_S10_M5 0
`define AXI_AR_LAYER_S10_M6 0
`define AXI_AR_LAYER_S10_M7 0
`define AXI_AR_LAYER_S10_M8 0
`define AXI_AR_LAYER_S10_M9 0
`define AXI_AR_LAYER_S10_M10 0
`define AXI_AR_LAYER_S10_M11 0
`define AXI_AR_LAYER_S10_M12 0
`define AXI_AR_LAYER_S10_M13 0
`define AXI_AR_LAYER_S10_M14 0
`define AXI_AR_LAYER_S10_M15 0
`define AXI_AR_LAYER_S10_M16 0
`define AXI_AW_LAYER_S10_M1 0
`define AXI_AW_LAYER_S10_M2 0
`define AXI_AW_LAYER_S10_M3 0
`define AXI_AW_LAYER_S10_M4 0
`define AXI_AW_LAYER_S10_M5 0
`define AXI_AW_LAYER_S10_M6 0
`define AXI_AW_LAYER_S10_M7 0
`define AXI_AW_LAYER_S10_M8 0
`define AXI_AW_LAYER_S10_M9 0
`define AXI_AW_LAYER_S10_M10 0
`define AXI_AW_LAYER_S10_M11 0
`define AXI_AW_LAYER_S10_M12 0
`define AXI_AW_LAYER_S10_M13 0
`define AXI_AW_LAYER_S10_M14 0
`define AXI_AW_LAYER_S10_M15 0
`define AXI_AW_LAYER_S10_M16 0
`define AXI_W_LAYER_S10_M1 0
`define AXI_W_LAYER_S10_M2 0
`define AXI_W_LAYER_S10_M3 0
`define AXI_W_LAYER_S10_M4 0
`define AXI_W_LAYER_S10_M5 0
`define AXI_W_LAYER_S10_M6 0
`define AXI_W_LAYER_S10_M7 0
`define AXI_W_LAYER_S10_M8 0
`define AXI_W_LAYER_S10_M9 0
`define AXI_W_LAYER_S10_M10 0
`define AXI_W_LAYER_S10_M11 0
`define AXI_W_LAYER_S10_M12 0
`define AXI_W_LAYER_S10_M13 0
`define AXI_W_LAYER_S10_M14 0
`define AXI_W_LAYER_S10_M15 0
`define AXI_W_LAYER_S10_M16 0
`define AXI_AR_LAYER_S11_M1 0
`define AXI_AR_LAYER_S11_M2 0
`define AXI_AR_LAYER_S11_M3 0
`define AXI_AR_LAYER_S11_M4 0
`define AXI_AR_LAYER_S11_M5 0
`define AXI_AR_LAYER_S11_M6 0
`define AXI_AR_LAYER_S11_M7 0
`define AXI_AR_LAYER_S11_M8 0
`define AXI_AR_LAYER_S11_M9 0
`define AXI_AR_LAYER_S11_M10 0
`define AXI_AR_LAYER_S11_M11 0
`define AXI_AR_LAYER_S11_M12 0
`define AXI_AR_LAYER_S11_M13 0
`define AXI_AR_LAYER_S11_M14 0
`define AXI_AR_LAYER_S11_M15 0
`define AXI_AR_LAYER_S11_M16 0
`define AXI_AW_LAYER_S11_M1 0
`define AXI_AW_LAYER_S11_M2 0
`define AXI_AW_LAYER_S11_M3 0
`define AXI_AW_LAYER_S11_M4 0
`define AXI_AW_LAYER_S11_M5 0
`define AXI_AW_LAYER_S11_M6 0
`define AXI_AW_LAYER_S11_M7 0
`define AXI_AW_LAYER_S11_M8 0
`define AXI_AW_LAYER_S11_M9 0
`define AXI_AW_LAYER_S11_M10 0
`define AXI_AW_LAYER_S11_M11 0
`define AXI_AW_LAYER_S11_M12 0
`define AXI_AW_LAYER_S11_M13 0
`define AXI_AW_LAYER_S11_M14 0
`define AXI_AW_LAYER_S11_M15 0
`define AXI_AW_LAYER_S11_M16 0
`define AXI_W_LAYER_S11_M1 0
`define AXI_W_LAYER_S11_M2 0
`define AXI_W_LAYER_S11_M3 0
`define AXI_W_LAYER_S11_M4 0
`define AXI_W_LAYER_S11_M5 0
`define AXI_W_LAYER_S11_M6 0
`define AXI_W_LAYER_S11_M7 0
`define AXI_W_LAYER_S11_M8 0
`define AXI_W_LAYER_S11_M9 0
`define AXI_W_LAYER_S11_M10 0
`define AXI_W_LAYER_S11_M11 0
`define AXI_W_LAYER_S11_M12 0
`define AXI_W_LAYER_S11_M13 0
`define AXI_W_LAYER_S11_M14 0
`define AXI_W_LAYER_S11_M15 0
`define AXI_W_LAYER_S11_M16 0
`define AXI_AR_LAYER_S12_M1 0
`define AXI_AR_LAYER_S12_M2 0
`define AXI_AR_LAYER_S12_M3 0
`define AXI_AR_LAYER_S12_M4 0
`define AXI_AR_LAYER_S12_M5 0
`define AXI_AR_LAYER_S12_M6 0
`define AXI_AR_LAYER_S12_M7 0
`define AXI_AR_LAYER_S12_M8 0
`define AXI_AR_LAYER_S12_M9 0
`define AXI_AR_LAYER_S12_M10 0
`define AXI_AR_LAYER_S12_M11 0
`define AXI_AR_LAYER_S12_M12 0
`define AXI_AR_LAYER_S12_M13 0
`define AXI_AR_LAYER_S12_M14 0
`define AXI_AR_LAYER_S12_M15 0
`define AXI_AR_LAYER_S12_M16 0
`define AXI_AW_LAYER_S12_M1 0
`define AXI_AW_LAYER_S12_M2 0
`define AXI_AW_LAYER_S12_M3 0
`define AXI_AW_LAYER_S12_M4 0
`define AXI_AW_LAYER_S12_M5 0
`define AXI_AW_LAYER_S12_M6 0
`define AXI_AW_LAYER_S12_M7 0
`define AXI_AW_LAYER_S12_M8 0
`define AXI_AW_LAYER_S12_M9 0
`define AXI_AW_LAYER_S12_M10 0
`define AXI_AW_LAYER_S12_M11 0
`define AXI_AW_LAYER_S12_M12 0
`define AXI_AW_LAYER_S12_M13 0
`define AXI_AW_LAYER_S12_M14 0
`define AXI_AW_LAYER_S12_M15 0
`define AXI_AW_LAYER_S12_M16 0
`define AXI_W_LAYER_S12_M1 0
`define AXI_W_LAYER_S12_M2 0
`define AXI_W_LAYER_S12_M3 0
`define AXI_W_LAYER_S12_M4 0
`define AXI_W_LAYER_S12_M5 0
`define AXI_W_LAYER_S12_M6 0
`define AXI_W_LAYER_S12_M7 0
`define AXI_W_LAYER_S12_M8 0
`define AXI_W_LAYER_S12_M9 0
`define AXI_W_LAYER_S12_M10 0
`define AXI_W_LAYER_S12_M11 0
`define AXI_W_LAYER_S12_M12 0
`define AXI_W_LAYER_S12_M13 0
`define AXI_W_LAYER_S12_M14 0
`define AXI_W_LAYER_S12_M15 0
`define AXI_W_LAYER_S12_M16 0
`define AXI_AR_LAYER_S13_M1 0
`define AXI_AR_LAYER_S13_M2 0
`define AXI_AR_LAYER_S13_M3 0
`define AXI_AR_LAYER_S13_M4 0
`define AXI_AR_LAYER_S13_M5 0
`define AXI_AR_LAYER_S13_M6 0
`define AXI_AR_LAYER_S13_M7 0
`define AXI_AR_LAYER_S13_M8 0
`define AXI_AR_LAYER_S13_M9 0
`define AXI_AR_LAYER_S13_M10 0
`define AXI_AR_LAYER_S13_M11 0
`define AXI_AR_LAYER_S13_M12 0
`define AXI_AR_LAYER_S13_M13 0
`define AXI_AR_LAYER_S13_M14 0
`define AXI_AR_LAYER_S13_M15 0
`define AXI_AR_LAYER_S13_M16 0
`define AXI_AW_LAYER_S13_M1 0
`define AXI_AW_LAYER_S13_M2 0
`define AXI_AW_LAYER_S13_M3 0
`define AXI_AW_LAYER_S13_M4 0
`define AXI_AW_LAYER_S13_M5 0
`define AXI_AW_LAYER_S13_M6 0
`define AXI_AW_LAYER_S13_M7 0
`define AXI_AW_LAYER_S13_M8 0
`define AXI_AW_LAYER_S13_M9 0
`define AXI_AW_LAYER_S13_M10 0
`define AXI_AW_LAYER_S13_M11 0
`define AXI_AW_LAYER_S13_M12 0
`define AXI_AW_LAYER_S13_M13 0
`define AXI_AW_LAYER_S13_M14 0
`define AXI_AW_LAYER_S13_M15 0
`define AXI_AW_LAYER_S13_M16 0
`define AXI_W_LAYER_S13_M1 0
`define AXI_W_LAYER_S13_M2 0
`define AXI_W_LAYER_S13_M3 0
`define AXI_W_LAYER_S13_M4 0
`define AXI_W_LAYER_S13_M5 0
`define AXI_W_LAYER_S13_M6 0
`define AXI_W_LAYER_S13_M7 0
`define AXI_W_LAYER_S13_M8 0
`define AXI_W_LAYER_S13_M9 0
`define AXI_W_LAYER_S13_M10 0
`define AXI_W_LAYER_S13_M11 0
`define AXI_W_LAYER_S13_M12 0
`define AXI_W_LAYER_S13_M13 0
`define AXI_W_LAYER_S13_M14 0
`define AXI_W_LAYER_S13_M15 0
`define AXI_W_LAYER_S13_M16 0
`define AXI_AR_LAYER_S14_M1 0
`define AXI_AR_LAYER_S14_M2 0
`define AXI_AR_LAYER_S14_M3 0
`define AXI_AR_LAYER_S14_M4 0
`define AXI_AR_LAYER_S14_M5 0
`define AXI_AR_LAYER_S14_M6 0
`define AXI_AR_LAYER_S14_M7 0
`define AXI_AR_LAYER_S14_M8 0
`define AXI_AR_LAYER_S14_M9 0
`define AXI_AR_LAYER_S14_M10 0
`define AXI_AR_LAYER_S14_M11 0
`define AXI_AR_LAYER_S14_M12 0
`define AXI_AR_LAYER_S14_M13 0
`define AXI_AR_LAYER_S14_M14 0
`define AXI_AR_LAYER_S14_M15 0
`define AXI_AR_LAYER_S14_M16 0
`define AXI_AW_LAYER_S14_M1 0
`define AXI_AW_LAYER_S14_M2 0
`define AXI_AW_LAYER_S14_M3 0
`define AXI_AW_LAYER_S14_M4 0
`define AXI_AW_LAYER_S14_M5 0
`define AXI_AW_LAYER_S14_M6 0
`define AXI_AW_LAYER_S14_M7 0
`define AXI_AW_LAYER_S14_M8 0
`define AXI_AW_LAYER_S14_M9 0
`define AXI_AW_LAYER_S14_M10 0
`define AXI_AW_LAYER_S14_M11 0
`define AXI_AW_LAYER_S14_M12 0
`define AXI_AW_LAYER_S14_M13 0
`define AXI_AW_LAYER_S14_M14 0
`define AXI_AW_LAYER_S14_M15 0
`define AXI_AW_LAYER_S14_M16 0
`define AXI_W_LAYER_S14_M1 0
`define AXI_W_LAYER_S14_M2 0
`define AXI_W_LAYER_S14_M3 0
`define AXI_W_LAYER_S14_M4 0
`define AXI_W_LAYER_S14_M5 0
`define AXI_W_LAYER_S14_M6 0
`define AXI_W_LAYER_S14_M7 0
`define AXI_W_LAYER_S14_M8 0
`define AXI_W_LAYER_S14_M9 0
`define AXI_W_LAYER_S14_M10 0
`define AXI_W_LAYER_S14_M11 0
`define AXI_W_LAYER_S14_M12 0
`define AXI_W_LAYER_S14_M13 0
`define AXI_W_LAYER_S14_M14 0
`define AXI_W_LAYER_S14_M15 0
`define AXI_W_LAYER_S14_M16 0
`define AXI_AR_LAYER_S15_M1 0
`define AXI_AR_LAYER_S15_M2 0
`define AXI_AR_LAYER_S15_M3 0
`define AXI_AR_LAYER_S15_M4 0
`define AXI_AR_LAYER_S15_M5 0
`define AXI_AR_LAYER_S15_M6 0
`define AXI_AR_LAYER_S15_M7 0
`define AXI_AR_LAYER_S15_M8 0
`define AXI_AR_LAYER_S15_M9 0
`define AXI_AR_LAYER_S15_M10 0
`define AXI_AR_LAYER_S15_M11 0
`define AXI_AR_LAYER_S15_M12 0
`define AXI_AR_LAYER_S15_M13 0
`define AXI_AR_LAYER_S15_M14 0
`define AXI_AR_LAYER_S15_M15 0
`define AXI_AR_LAYER_S15_M16 0
`define AXI_AW_LAYER_S15_M1 0
`define AXI_AW_LAYER_S15_M2 0
`define AXI_AW_LAYER_S15_M3 0
`define AXI_AW_LAYER_S15_M4 0
`define AXI_AW_LAYER_S15_M5 0
`define AXI_AW_LAYER_S15_M6 0
`define AXI_AW_LAYER_S15_M7 0
`define AXI_AW_LAYER_S15_M8 0
`define AXI_AW_LAYER_S15_M9 0
`define AXI_AW_LAYER_S15_M10 0
`define AXI_AW_LAYER_S15_M11 0
`define AXI_AW_LAYER_S15_M12 0
`define AXI_AW_LAYER_S15_M13 0
`define AXI_AW_LAYER_S15_M14 0
`define AXI_AW_LAYER_S15_M15 0
`define AXI_AW_LAYER_S15_M16 0
`define AXI_W_LAYER_S15_M1 0
`define AXI_W_LAYER_S15_M2 0
`define AXI_W_LAYER_S15_M3 0
`define AXI_W_LAYER_S15_M4 0
`define AXI_W_LAYER_S15_M5 0
`define AXI_W_LAYER_S15_M6 0
`define AXI_W_LAYER_S15_M7 0
`define AXI_W_LAYER_S15_M8 0
`define AXI_W_LAYER_S15_M9 0
`define AXI_W_LAYER_S15_M10 0
`define AXI_W_LAYER_S15_M11 0
`define AXI_W_LAYER_S15_M12 0
`define AXI_W_LAYER_S15_M13 0
`define AXI_W_LAYER_S15_M14 0
`define AXI_W_LAYER_S15_M15 0
`define AXI_W_LAYER_S15_M16 0
`define AXI_AR_LAYER_S16_M1 0
`define AXI_AR_LAYER_S16_M2 0
`define AXI_AR_LAYER_S16_M3 0
`define AXI_AR_LAYER_S16_M4 0
`define AXI_AR_LAYER_S16_M5 0
`define AXI_AR_LAYER_S16_M6 0
`define AXI_AR_LAYER_S16_M7 0
`define AXI_AR_LAYER_S16_M8 0
`define AXI_AR_LAYER_S16_M9 0
`define AXI_AR_LAYER_S16_M10 0
`define AXI_AR_LAYER_S16_M11 0
`define AXI_AR_LAYER_S16_M12 0
`define AXI_AR_LAYER_S16_M13 0
`define AXI_AR_LAYER_S16_M14 0
`define AXI_AR_LAYER_S16_M15 0
`define AXI_AR_LAYER_S16_M16 0
`define AXI_AW_LAYER_S16_M1 0
`define AXI_AW_LAYER_S16_M2 0
`define AXI_AW_LAYER_S16_M3 0
`define AXI_AW_LAYER_S16_M4 0
`define AXI_AW_LAYER_S16_M5 0
`define AXI_AW_LAYER_S16_M6 0
`define AXI_AW_LAYER_S16_M7 0
`define AXI_AW_LAYER_S16_M8 0
`define AXI_AW_LAYER_S16_M9 0
`define AXI_AW_LAYER_S16_M10 0
`define AXI_AW_LAYER_S16_M11 0
`define AXI_AW_LAYER_S16_M12 0
`define AXI_AW_LAYER_S16_M13 0
`define AXI_AW_LAYER_S16_M14 0
`define AXI_AW_LAYER_S16_M15 0
`define AXI_AW_LAYER_S16_M16 0
`define AXI_W_LAYER_S16_M1 0
`define AXI_W_LAYER_S16_M2 0
`define AXI_W_LAYER_S16_M3 0
`define AXI_W_LAYER_S16_M4 0
`define AXI_W_LAYER_S16_M5 0
`define AXI_W_LAYER_S16_M6 0
`define AXI_W_LAYER_S16_M7 0
`define AXI_W_LAYER_S16_M8 0
`define AXI_W_LAYER_S16_M9 0
`define AXI_W_LAYER_S16_M10 0
`define AXI_W_LAYER_S16_M11 0
`define AXI_W_LAYER_S16_M12 0
`define AXI_W_LAYER_S16_M13 0
`define AXI_W_LAYER_S16_M14 0
`define AXI_W_LAYER_S16_M15 0
`define AXI_W_LAYER_S16_M16 0
`define AXI_ALL_R_LAYER_SHARED 0
`define AXI_R_LAYER_M1_S0 0
`define AXI_R_LAYER_M1_S1 0
`define AXI_R_LAYER_M1_S2 0
`define AXI_R_LAYER_M1_S3 0
`define AXI_R_LAYER_M1_S4 0
`define AXI_R_LAYER_M1_S5 0
`define AXI_R_LAYER_M1_S6 0
`define AXI_R_LAYER_M1_S7 0
`define AXI_R_LAYER_M1_S8 0
`define AXI_R_LAYER_M1_S9 0
`define AXI_R_LAYER_M1_S10 0
`define AXI_R_LAYER_M1_S11 0
`define AXI_R_LAYER_M1_S12 0
`define AXI_R_LAYER_M1_S13 0
`define AXI_R_LAYER_M1_S14 0
`define AXI_R_LAYER_M1_S15 0
`define AXI_R_LAYER_M1_S16 0
`define AXI_ALL_B_LAYER_SHARED 0
`define AXI_B_LAYER_M1_S0 0
`define AXI_B_LAYER_M1_S1 0
`define AXI_B_LAYER_M1_S2 0
`define AXI_B_LAYER_M1_S3 0
`define AXI_B_LAYER_M1_S4 0
`define AXI_B_LAYER_M1_S5 0
`define AXI_B_LAYER_M1_S6 0
`define AXI_B_LAYER_M1_S7 0
`define AXI_B_LAYER_M1_S8 0
`define AXI_B_LAYER_M1_S9 0
`define AXI_B_LAYER_M1_S10 0
`define AXI_B_LAYER_M1_S11 0
`define AXI_B_LAYER_M1_S12 0
`define AXI_B_LAYER_M1_S13 0
`define AXI_B_LAYER_M1_S14 0
`define AXI_B_LAYER_M1_S15 0
`define AXI_B_LAYER_M1_S16 0
`define AXI_R_LAYER_M2_S0 0
`define AXI_R_LAYER_M2_S1 0
`define AXI_R_LAYER_M2_S2 0
`define AXI_R_LAYER_M2_S3 0
`define AXI_R_LAYER_M2_S4 0
`define AXI_R_LAYER_M2_S5 0
`define AXI_R_LAYER_M2_S6 0
`define AXI_R_LAYER_M2_S7 0
`define AXI_R_LAYER_M2_S8 0
`define AXI_R_LAYER_M2_S9 0
`define AXI_R_LAYER_M2_S10 0
`define AXI_R_LAYER_M2_S11 0
`define AXI_R_LAYER_M2_S12 0
`define AXI_R_LAYER_M2_S13 0
`define AXI_R_LAYER_M2_S14 0
`define AXI_R_LAYER_M2_S15 0
`define AXI_R_LAYER_M2_S16 0
`define AXI_B_LAYER_M2_S0 0
`define AXI_B_LAYER_M2_S1 0
`define AXI_B_LAYER_M2_S2 0
`define AXI_B_LAYER_M2_S3 0
`define AXI_B_LAYER_M2_S4 0
`define AXI_B_LAYER_M2_S5 0
`define AXI_B_LAYER_M2_S6 0
`define AXI_B_LAYER_M2_S7 0
`define AXI_B_LAYER_M2_S8 0
`define AXI_B_LAYER_M2_S9 0
`define AXI_B_LAYER_M2_S10 0
`define AXI_B_LAYER_M2_S11 0
`define AXI_B_LAYER_M2_S12 0
`define AXI_B_LAYER_M2_S13 0
`define AXI_B_LAYER_M2_S14 0
`define AXI_B_LAYER_M2_S15 0
`define AXI_B_LAYER_M2_S16 0
`define AXI_R_LAYER_M3_S0 0
`define AXI_R_LAYER_M3_S1 0
`define AXI_R_LAYER_M3_S2 0
`define AXI_R_LAYER_M3_S3 0
`define AXI_R_LAYER_M3_S4 0
`define AXI_R_LAYER_M3_S5 0
`define AXI_R_LAYER_M3_S6 0
`define AXI_R_LAYER_M3_S7 0
`define AXI_R_LAYER_M3_S8 0
`define AXI_R_LAYER_M3_S9 0
`define AXI_R_LAYER_M3_S10 0
`define AXI_R_LAYER_M3_S11 0
`define AXI_R_LAYER_M3_S12 0
`define AXI_R_LAYER_M3_S13 0
`define AXI_R_LAYER_M3_S14 0
`define AXI_R_LAYER_M3_S15 0
`define AXI_R_LAYER_M3_S16 0
`define AXI_B_LAYER_M3_S0 0
`define AXI_B_LAYER_M3_S1 0
`define AXI_B_LAYER_M3_S2 0
`define AXI_B_LAYER_M3_S3 0
`define AXI_B_LAYER_M3_S4 0
`define AXI_B_LAYER_M3_S5 0
`define AXI_B_LAYER_M3_S6 0
`define AXI_B_LAYER_M3_S7 0
`define AXI_B_LAYER_M3_S8 0
`define AXI_B_LAYER_M3_S9 0
`define AXI_B_LAYER_M3_S10 0
`define AXI_B_LAYER_M3_S11 0
`define AXI_B_LAYER_M3_S12 0
`define AXI_B_LAYER_M3_S13 0
`define AXI_B_LAYER_M3_S14 0
`define AXI_B_LAYER_M3_S15 0
`define AXI_B_LAYER_M3_S16 0
`define AXI_R_LAYER_M4_S0 0
`define AXI_R_LAYER_M4_S1 0
`define AXI_R_LAYER_M4_S2 0
`define AXI_R_LAYER_M4_S3 0
`define AXI_R_LAYER_M4_S4 0
`define AXI_R_LAYER_M4_S5 0
`define AXI_R_LAYER_M4_S6 0
`define AXI_R_LAYER_M4_S7 0
`define AXI_R_LAYER_M4_S8 0
`define AXI_R_LAYER_M4_S9 0
`define AXI_R_LAYER_M4_S10 0
`define AXI_R_LAYER_M4_S11 0
`define AXI_R_LAYER_M4_S12 0
`define AXI_R_LAYER_M4_S13 0
`define AXI_R_LAYER_M4_S14 0
`define AXI_R_LAYER_M4_S15 0
`define AXI_R_LAYER_M4_S16 0
`define AXI_B_LAYER_M4_S0 0
`define AXI_B_LAYER_M4_S1 0
`define AXI_B_LAYER_M4_S2 0
`define AXI_B_LAYER_M4_S3 0
`define AXI_B_LAYER_M4_S4 0
`define AXI_B_LAYER_M4_S5 0
`define AXI_B_LAYER_M4_S6 0
`define AXI_B_LAYER_M4_S7 0
`define AXI_B_LAYER_M4_S8 0
`define AXI_B_LAYER_M4_S9 0
`define AXI_B_LAYER_M4_S10 0
`define AXI_B_LAYER_M4_S11 0
`define AXI_B_LAYER_M4_S12 0
`define AXI_B_LAYER_M4_S13 0
`define AXI_B_LAYER_M4_S14 0
`define AXI_B_LAYER_M4_S15 0
`define AXI_B_LAYER_M4_S16 0
`define AXI_R_LAYER_M5_S0 0
`define AXI_R_LAYER_M5_S1 0
`define AXI_R_LAYER_M5_S2 0
`define AXI_R_LAYER_M5_S3 0
`define AXI_R_LAYER_M5_S4 0
`define AXI_R_LAYER_M5_S5 0
`define AXI_R_LAYER_M5_S6 0
`define AXI_R_LAYER_M5_S7 0
`define AXI_R_LAYER_M5_S8 0
`define AXI_R_LAYER_M5_S9 0
`define AXI_R_LAYER_M5_S10 0
`define AXI_R_LAYER_M5_S11 0
`define AXI_R_LAYER_M5_S12 0
`define AXI_R_LAYER_M5_S13 0
`define AXI_R_LAYER_M5_S14 0
`define AXI_R_LAYER_M5_S15 0
`define AXI_R_LAYER_M5_S16 0
`define AXI_B_LAYER_M5_S0 0
`define AXI_B_LAYER_M5_S1 0
`define AXI_B_LAYER_M5_S2 0
`define AXI_B_LAYER_M5_S3 0
`define AXI_B_LAYER_M5_S4 0
`define AXI_B_LAYER_M5_S5 0
`define AXI_B_LAYER_M5_S6 0
`define AXI_B_LAYER_M5_S7 0
`define AXI_B_LAYER_M5_S8 0
`define AXI_B_LAYER_M5_S9 0
`define AXI_B_LAYER_M5_S10 0
`define AXI_B_LAYER_M5_S11 0
`define AXI_B_LAYER_M5_S12 0
`define AXI_B_LAYER_M5_S13 0
`define AXI_B_LAYER_M5_S14 0
`define AXI_B_LAYER_M5_S15 0
`define AXI_B_LAYER_M5_S16 0
`define AXI_R_LAYER_M6_S0 0
`define AXI_R_LAYER_M6_S1 0
`define AXI_R_LAYER_M6_S2 0
`define AXI_R_LAYER_M6_S3 0
`define AXI_R_LAYER_M6_S4 0
`define AXI_R_LAYER_M6_S5 0
`define AXI_R_LAYER_M6_S6 0
`define AXI_R_LAYER_M6_S7 0
`define AXI_R_LAYER_M6_S8 0
`define AXI_R_LAYER_M6_S9 0
`define AXI_R_LAYER_M6_S10 0
`define AXI_R_LAYER_M6_S11 0
`define AXI_R_LAYER_M6_S12 0
`define AXI_R_LAYER_M6_S13 0
`define AXI_R_LAYER_M6_S14 0
`define AXI_R_LAYER_M6_S15 0
`define AXI_R_LAYER_M6_S16 0
`define AXI_B_LAYER_M6_S0 0
`define AXI_B_LAYER_M6_S1 0
`define AXI_B_LAYER_M6_S2 0
`define AXI_B_LAYER_M6_S3 0
`define AXI_B_LAYER_M6_S4 0
`define AXI_B_LAYER_M6_S5 0
`define AXI_B_LAYER_M6_S6 0
`define AXI_B_LAYER_M6_S7 0
`define AXI_B_LAYER_M6_S8 0
`define AXI_B_LAYER_M6_S9 0
`define AXI_B_LAYER_M6_S10 0
`define AXI_B_LAYER_M6_S11 0
`define AXI_B_LAYER_M6_S12 0
`define AXI_B_LAYER_M6_S13 0
`define AXI_B_LAYER_M6_S14 0
`define AXI_B_LAYER_M6_S15 0
`define AXI_B_LAYER_M6_S16 0
`define AXI_R_LAYER_M7_S0 0
`define AXI_R_LAYER_M7_S1 0
`define AXI_R_LAYER_M7_S2 0
`define AXI_R_LAYER_M7_S3 0
`define AXI_R_LAYER_M7_S4 0
`define AXI_R_LAYER_M7_S5 0
`define AXI_R_LAYER_M7_S6 0
`define AXI_R_LAYER_M7_S7 0
`define AXI_R_LAYER_M7_S8 0
`define AXI_R_LAYER_M7_S9 0
`define AXI_R_LAYER_M7_S10 0
`define AXI_R_LAYER_M7_S11 0
`define AXI_R_LAYER_M7_S12 0
`define AXI_R_LAYER_M7_S13 0
`define AXI_R_LAYER_M7_S14 0
`define AXI_R_LAYER_M7_S15 0
`define AXI_R_LAYER_M7_S16 0
`define AXI_B_LAYER_M7_S0 0
`define AXI_B_LAYER_M7_S1 0
`define AXI_B_LAYER_M7_S2 0
`define AXI_B_LAYER_M7_S3 0
`define AXI_B_LAYER_M7_S4 0
`define AXI_B_LAYER_M7_S5 0
`define AXI_B_LAYER_M7_S6 0
`define AXI_B_LAYER_M7_S7 0
`define AXI_B_LAYER_M7_S8 0
`define AXI_B_LAYER_M7_S9 0
`define AXI_B_LAYER_M7_S10 0
`define AXI_B_LAYER_M7_S11 0
`define AXI_B_LAYER_M7_S12 0
`define AXI_B_LAYER_M7_S13 0
`define AXI_B_LAYER_M7_S14 0
`define AXI_B_LAYER_M7_S15 0
`define AXI_B_LAYER_M7_S16 0
`define AXI_R_LAYER_M8_S0 0
`define AXI_R_LAYER_M8_S1 0
`define AXI_R_LAYER_M8_S2 0
`define AXI_R_LAYER_M8_S3 0
`define AXI_R_LAYER_M8_S4 0
`define AXI_R_LAYER_M8_S5 0
`define AXI_R_LAYER_M8_S6 0
`define AXI_R_LAYER_M8_S7 0
`define AXI_R_LAYER_M8_S8 0
`define AXI_R_LAYER_M8_S9 0
`define AXI_R_LAYER_M8_S10 0
`define AXI_R_LAYER_M8_S11 0
`define AXI_R_LAYER_M8_S12 0
`define AXI_R_LAYER_M8_S13 0
`define AXI_R_LAYER_M8_S14 0
`define AXI_R_LAYER_M8_S15 0
`define AXI_R_LAYER_M8_S16 0
`define AXI_B_LAYER_M8_S0 0
`define AXI_B_LAYER_M8_S1 0
`define AXI_B_LAYER_M8_S2 0
`define AXI_B_LAYER_M8_S3 0
`define AXI_B_LAYER_M8_S4 0
`define AXI_B_LAYER_M8_S5 0
`define AXI_B_LAYER_M8_S6 0
`define AXI_B_LAYER_M8_S7 0
`define AXI_B_LAYER_M8_S8 0
`define AXI_B_LAYER_M8_S9 0
`define AXI_B_LAYER_M8_S10 0
`define AXI_B_LAYER_M8_S11 0
`define AXI_B_LAYER_M8_S12 0
`define AXI_B_LAYER_M8_S13 0
`define AXI_B_LAYER_M8_S14 0
`define AXI_B_LAYER_M8_S15 0
`define AXI_B_LAYER_M8_S16 0
`define AXI_R_LAYER_M9_S0 0
`define AXI_R_LAYER_M9_S1 0
`define AXI_R_LAYER_M9_S2 0
`define AXI_R_LAYER_M9_S3 0
`define AXI_R_LAYER_M9_S4 0
`define AXI_R_LAYER_M9_S5 0
`define AXI_R_LAYER_M9_S6 0
`define AXI_R_LAYER_M9_S7 0
`define AXI_R_LAYER_M9_S8 0
`define AXI_R_LAYER_M9_S9 0
`define AXI_R_LAYER_M9_S10 0
`define AXI_R_LAYER_M9_S11 0
`define AXI_R_LAYER_M9_S12 0
`define AXI_R_LAYER_M9_S13 0
`define AXI_R_LAYER_M9_S14 0
`define AXI_R_LAYER_M9_S15 0
`define AXI_R_LAYER_M9_S16 0
`define AXI_B_LAYER_M9_S0 0
`define AXI_B_LAYER_M9_S1 0
`define AXI_B_LAYER_M9_S2 0
`define AXI_B_LAYER_M9_S3 0
`define AXI_B_LAYER_M9_S4 0
`define AXI_B_LAYER_M9_S5 0
`define AXI_B_LAYER_M9_S6 0
`define AXI_B_LAYER_M9_S7 0
`define AXI_B_LAYER_M9_S8 0
`define AXI_B_LAYER_M9_S9 0
`define AXI_B_LAYER_M9_S10 0
`define AXI_B_LAYER_M9_S11 0
`define AXI_B_LAYER_M9_S12 0
`define AXI_B_LAYER_M9_S13 0
`define AXI_B_LAYER_M9_S14 0
`define AXI_B_LAYER_M9_S15 0
`define AXI_B_LAYER_M9_S16 0
`define AXI_R_LAYER_M10_S0 0
`define AXI_R_LAYER_M10_S1 0
`define AXI_R_LAYER_M10_S2 0
`define AXI_R_LAYER_M10_S3 0
`define AXI_R_LAYER_M10_S4 0
`define AXI_R_LAYER_M10_S5 0
`define AXI_R_LAYER_M10_S6 0
`define AXI_R_LAYER_M10_S7 0
`define AXI_R_LAYER_M10_S8 0
`define AXI_R_LAYER_M10_S9 0
`define AXI_R_LAYER_M10_S10 0
`define AXI_R_LAYER_M10_S11 0
`define AXI_R_LAYER_M10_S12 0
`define AXI_R_LAYER_M10_S13 0
`define AXI_R_LAYER_M10_S14 0
`define AXI_R_LAYER_M10_S15 0
`define AXI_R_LAYER_M10_S16 0
`define AXI_B_LAYER_M10_S0 0
`define AXI_B_LAYER_M10_S1 0
`define AXI_B_LAYER_M10_S2 0
`define AXI_B_LAYER_M10_S3 0
`define AXI_B_LAYER_M10_S4 0
`define AXI_B_LAYER_M10_S5 0
`define AXI_B_LAYER_M10_S6 0
`define AXI_B_LAYER_M10_S7 0
`define AXI_B_LAYER_M10_S8 0
`define AXI_B_LAYER_M10_S9 0
`define AXI_B_LAYER_M10_S10 0
`define AXI_B_LAYER_M10_S11 0
`define AXI_B_LAYER_M10_S12 0
`define AXI_B_LAYER_M10_S13 0
`define AXI_B_LAYER_M10_S14 0
`define AXI_B_LAYER_M10_S15 0
`define AXI_B_LAYER_M10_S16 0
`define AXI_R_LAYER_M11_S0 0
`define AXI_R_LAYER_M11_S1 0
`define AXI_R_LAYER_M11_S2 0
`define AXI_R_LAYER_M11_S3 0
`define AXI_R_LAYER_M11_S4 0
`define AXI_R_LAYER_M11_S5 0
`define AXI_R_LAYER_M11_S6 0
`define AXI_R_LAYER_M11_S7 0
`define AXI_R_LAYER_M11_S8 0
`define AXI_R_LAYER_M11_S9 0
`define AXI_R_LAYER_M11_S10 0
`define AXI_R_LAYER_M11_S11 0
`define AXI_R_LAYER_M11_S12 0
`define AXI_R_LAYER_M11_S13 0
`define AXI_R_LAYER_M11_S14 0
`define AXI_R_LAYER_M11_S15 0
`define AXI_R_LAYER_M11_S16 0
`define AXI_B_LAYER_M11_S0 0
`define AXI_B_LAYER_M11_S1 0
`define AXI_B_LAYER_M11_S2 0
`define AXI_B_LAYER_M11_S3 0
`define AXI_B_LAYER_M11_S4 0
`define AXI_B_LAYER_M11_S5 0
`define AXI_B_LAYER_M11_S6 0
`define AXI_B_LAYER_M11_S7 0
`define AXI_B_LAYER_M11_S8 0
`define AXI_B_LAYER_M11_S9 0
`define AXI_B_LAYER_M11_S10 0
`define AXI_B_LAYER_M11_S11 0
`define AXI_B_LAYER_M11_S12 0
`define AXI_B_LAYER_M11_S13 0
`define AXI_B_LAYER_M11_S14 0
`define AXI_B_LAYER_M11_S15 0
`define AXI_B_LAYER_M11_S16 0
`define AXI_R_LAYER_M12_S0 0
`define AXI_R_LAYER_M12_S1 0
`define AXI_R_LAYER_M12_S2 0
`define AXI_R_LAYER_M12_S3 0
`define AXI_R_LAYER_M12_S4 0
`define AXI_R_LAYER_M12_S5 0
`define AXI_R_LAYER_M12_S6 0
`define AXI_R_LAYER_M12_S7 0
`define AXI_R_LAYER_M12_S8 0
`define AXI_R_LAYER_M12_S9 0
`define AXI_R_LAYER_M12_S10 0
`define AXI_R_LAYER_M12_S11 0
`define AXI_R_LAYER_M12_S12 0
`define AXI_R_LAYER_M12_S13 0
`define AXI_R_LAYER_M12_S14 0
`define AXI_R_LAYER_M12_S15 0
`define AXI_R_LAYER_M12_S16 0
`define AXI_B_LAYER_M12_S0 0
`define AXI_B_LAYER_M12_S1 0
`define AXI_B_LAYER_M12_S2 0
`define AXI_B_LAYER_M12_S3 0
`define AXI_B_LAYER_M12_S4 0
`define AXI_B_LAYER_M12_S5 0
`define AXI_B_LAYER_M12_S6 0
`define AXI_B_LAYER_M12_S7 0
`define AXI_B_LAYER_M12_S8 0
`define AXI_B_LAYER_M12_S9 0
`define AXI_B_LAYER_M12_S10 0
`define AXI_B_LAYER_M12_S11 0
`define AXI_B_LAYER_M12_S12 0
`define AXI_B_LAYER_M12_S13 0
`define AXI_B_LAYER_M12_S14 0
`define AXI_B_LAYER_M12_S15 0
`define AXI_B_LAYER_M12_S16 0
`define AXI_R_LAYER_M13_S0 0
`define AXI_R_LAYER_M13_S1 0
`define AXI_R_LAYER_M13_S2 0
`define AXI_R_LAYER_M13_S3 0
`define AXI_R_LAYER_M13_S4 0
`define AXI_R_LAYER_M13_S5 0
`define AXI_R_LAYER_M13_S6 0
`define AXI_R_LAYER_M13_S7 0
`define AXI_R_LAYER_M13_S8 0
`define AXI_R_LAYER_M13_S9 0
`define AXI_R_LAYER_M13_S10 0
`define AXI_R_LAYER_M13_S11 0
`define AXI_R_LAYER_M13_S12 0
`define AXI_R_LAYER_M13_S13 0
`define AXI_R_LAYER_M13_S14 0
`define AXI_R_LAYER_M13_S15 0
`define AXI_R_LAYER_M13_S16 0
`define AXI_B_LAYER_M13_S0 0
`define AXI_B_LAYER_M13_S1 0
`define AXI_B_LAYER_M13_S2 0
`define AXI_B_LAYER_M13_S3 0
`define AXI_B_LAYER_M13_S4 0
`define AXI_B_LAYER_M13_S5 0
`define AXI_B_LAYER_M13_S6 0
`define AXI_B_LAYER_M13_S7 0
`define AXI_B_LAYER_M13_S8 0
`define AXI_B_LAYER_M13_S9 0
`define AXI_B_LAYER_M13_S10 0
`define AXI_B_LAYER_M13_S11 0
`define AXI_B_LAYER_M13_S12 0
`define AXI_B_LAYER_M13_S13 0
`define AXI_B_LAYER_M13_S14 0
`define AXI_B_LAYER_M13_S15 0
`define AXI_B_LAYER_M13_S16 0
`define AXI_R_LAYER_M14_S0 0
`define AXI_R_LAYER_M14_S1 0
`define AXI_R_LAYER_M14_S2 0
`define AXI_R_LAYER_M14_S3 0
`define AXI_R_LAYER_M14_S4 0
`define AXI_R_LAYER_M14_S5 0
`define AXI_R_LAYER_M14_S6 0
`define AXI_R_LAYER_M14_S7 0
`define AXI_R_LAYER_M14_S8 0
`define AXI_R_LAYER_M14_S9 0
`define AXI_R_LAYER_M14_S10 0
`define AXI_R_LAYER_M14_S11 0
`define AXI_R_LAYER_M14_S12 0
`define AXI_R_LAYER_M14_S13 0
`define AXI_R_LAYER_M14_S14 0
`define AXI_R_LAYER_M14_S15 0
`define AXI_R_LAYER_M14_S16 0
`define AXI_B_LAYER_M14_S0 0
`define AXI_B_LAYER_M14_S1 0
`define AXI_B_LAYER_M14_S2 0
`define AXI_B_LAYER_M14_S3 0
`define AXI_B_LAYER_M14_S4 0
`define AXI_B_LAYER_M14_S5 0
`define AXI_B_LAYER_M14_S6 0
`define AXI_B_LAYER_M14_S7 0
`define AXI_B_LAYER_M14_S8 0
`define AXI_B_LAYER_M14_S9 0
`define AXI_B_LAYER_M14_S10 0
`define AXI_B_LAYER_M14_S11 0
`define AXI_B_LAYER_M14_S12 0
`define AXI_B_LAYER_M14_S13 0
`define AXI_B_LAYER_M14_S14 0
`define AXI_B_LAYER_M14_S15 0
`define AXI_B_LAYER_M14_S16 0
`define AXI_R_LAYER_M15_S0 0
`define AXI_R_LAYER_M15_S1 0
`define AXI_R_LAYER_M15_S2 0
`define AXI_R_LAYER_M15_S3 0
`define AXI_R_LAYER_M15_S4 0
`define AXI_R_LAYER_M15_S5 0
`define AXI_R_LAYER_M15_S6 0
`define AXI_R_LAYER_M15_S7 0
`define AXI_R_LAYER_M15_S8 0
`define AXI_R_LAYER_M15_S9 0
`define AXI_R_LAYER_M15_S10 0
`define AXI_R_LAYER_M15_S11 0
`define AXI_R_LAYER_M15_S12 0
`define AXI_R_LAYER_M15_S13 0
`define AXI_R_LAYER_M15_S14 0
`define AXI_R_LAYER_M15_S15 0
`define AXI_R_LAYER_M15_S16 0
`define AXI_B_LAYER_M15_S0 0
`define AXI_B_LAYER_M15_S1 0
`define AXI_B_LAYER_M15_S2 0
`define AXI_B_LAYER_M15_S3 0
`define AXI_B_LAYER_M15_S4 0
`define AXI_B_LAYER_M15_S5 0
`define AXI_B_LAYER_M15_S6 0
`define AXI_B_LAYER_M15_S7 0
`define AXI_B_LAYER_M15_S8 0
`define AXI_B_LAYER_M15_S9 0
`define AXI_B_LAYER_M15_S10 0
`define AXI_B_LAYER_M15_S11 0
`define AXI_B_LAYER_M15_S12 0
`define AXI_B_LAYER_M15_S13 0
`define AXI_B_LAYER_M15_S14 0
`define AXI_B_LAYER_M15_S15 0
`define AXI_B_LAYER_M15_S16 0
`define AXI_R_LAYER_M16_S0 0
`define AXI_R_LAYER_M16_S1 0
`define AXI_R_LAYER_M16_S2 0
`define AXI_R_LAYER_M16_S3 0
`define AXI_R_LAYER_M16_S4 0
`define AXI_R_LAYER_M16_S5 0
`define AXI_R_LAYER_M16_S6 0
`define AXI_R_LAYER_M16_S7 0
`define AXI_R_LAYER_M16_S8 0
`define AXI_R_LAYER_M16_S9 0
`define AXI_R_LAYER_M16_S10 0
`define AXI_R_LAYER_M16_S11 0
`define AXI_R_LAYER_M16_S12 0
`define AXI_R_LAYER_M16_S13 0
`define AXI_R_LAYER_M16_S14 0
`define AXI_R_LAYER_M16_S15 0
`define AXI_R_LAYER_M16_S16 0
`define AXI_B_LAYER_M16_S0 0
`define AXI_B_LAYER_M16_S1 0
`define AXI_B_LAYER_M16_S2 0
`define AXI_B_LAYER_M16_S3 0
`define AXI_B_LAYER_M16_S4 0
`define AXI_B_LAYER_M16_S5 0
`define AXI_B_LAYER_M16_S6 0
`define AXI_B_LAYER_M16_S7 0
`define AXI_B_LAYER_M16_S8 0
`define AXI_B_LAYER_M16_S9 0
`define AXI_B_LAYER_M16_S10 0
`define AXI_B_LAYER_M16_S11 0
`define AXI_B_LAYER_M16_S12 0
`define AXI_B_LAYER_M16_S13 0
`define AXI_B_LAYER_M16_S14 0
`define AXI_B_LAYER_M16_S15 0
`define AXI_B_LAYER_M16_S16 0
`define AXI_AR_HAS_SHARED_LAYER 0
`define AXI_AW_HAS_SHARED_LAYER 0
`define AXI_W_HAS_SHARED_LAYER 0
`define AXI_R_HAS_SHARED_LAYER 0
`define AXI_B_HAS_SHARED_LAYER 0
`define AXI_AR_SHARED_LAYER_NM 1
`define AXI_LOG2_AR_SHARED_LAYER_NM 1
`define AXI_LOG2_AR_SHARED_LAYER_NMP1 1
`define AXI_AR_SHARED_LAYER_NS 1
`define AXI_AR_SHARED_LAYER_NS_R0 0
`define AXI_LOG2_AR_SHARED_LAYER_NS 1
`define AXI_LOG2_AR_SHARED_LAYER_NSP1 1
`define AXI_AW_SHARED_LAYER_NM 1
`define AXI_LOG2_AW_SHARED_LAYER_NM 1
`define AXI_LOG2_AW_SHARED_LAYER_NMP1 1
`define AXI_AW_SHARED_LAYER_NS 1
`define AXI_AW_SHARED_LAYER_NS_R0 0
`define AXI_LOG2_AW_SHARED_LAYER_NS 1
`define AXI_LOG2_AW_SHARED_LAYER_NSP1 1
`define AXI_W_SHARED_LAYER_NM 1
`define AXI_LOG2_W_SHARED_LAYER_NM 1
`define AXI_LOG2_W_SHARED_LAYER_NMP1 1
`define AXI_W_SHARED_LAYER_NS 1
`define AXI_W_SHARED_LAYER_NS_R0 0
`define AXI_LOG2_W_SHARED_LAYER_NS 1
`define AXI_LOG2_W_SHARED_LAYER_NSP1 1
`define AXI_R_SHARED_LAYER_NM 1
`define AXI_R_SHARED_LAYER_NM_R0 0
`define AXI_LOG2_R_SHARED_LAYER_NM 1
`define AXI_LOG2_R_SHARED_LAYER_NMP1 1
`define AXI_R_SHARED_LAYER_NS 1
`define AXI_LOG2_R_SHARED_LAYER_NS 1
`define AXI_LOG2_R_SHARED_LAYER_NSP1 1
`define AXI_B_SHARED_LAYER_NM 1
`define AXI_B_SHARED_LAYER_NM_R0 0
`define AXI_LOG2_B_SHARED_LAYER_NM 1
`define AXI_LOG2_B_SHARED_LAYER_NMP1 1
`define AXI_B_SHARED_LAYER_NS 1
`define AXI_LOG2_B_SHARED_LAYER_NS 1
`define AXI_LOG2_B_SHARED_LAYER_NSP1 1
`define AXI_AR_S0_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AR_S0_NMV 2
`define AXI_AR_S0_NMV_LOG2 1
`define AXI_AR_S0_NMV_P1_LOG2 2
`define AXI_AW_S0_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AW_S0_NMV 2
`define AXI_AW_S0_NMV_LOG2 1
`define AXI_AW_S0_NMV_P1_LOG2 2
`define AXI_W_S0_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_W_S0_NMV 2
`define AXI_W_S0_NMV_LOG2 1
`define AXI_W_S0_NMV_P1_LOG2 2
`define AXI_AR_S1_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AR_S1_NMV 2
`define AXI_AR_S1_NMV_LOG2 1
`define AXI_AR_S1_NMV_P1_LOG2 2
`define AXI_AW_S1_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AW_S1_NMV 2
`define AXI_AW_S1_NMV_LOG2 1
`define AXI_AW_S1_NMV_P1_LOG2 2
`define AXI_W_S1_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_W_S1_NMV 2
`define AXI_W_S1_NMV_LOG2 1
`define AXI_W_S1_NMV_P1_LOG2 2
`define AXI_AR_S2_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AR_S2_NMV 2
`define AXI_AR_S2_NMV_LOG2 1
`define AXI_AR_S2_NMV_P1_LOG2 2
`define AXI_AW_S2_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AW_S2_NMV 2
`define AXI_AW_S2_NMV_LOG2 1
`define AXI_AW_S2_NMV_P1_LOG2 2
`define AXI_W_S2_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_W_S2_NMV 2
`define AXI_W_S2_NMV_LOG2 1
`define AXI_W_S2_NMV_P1_LOG2 2
`define AXI_AR_S3_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AR_S3_NMV 2
`define AXI_AR_S3_NMV_LOG2 1
`define AXI_AR_S3_NMV_P1_LOG2 2
`define AXI_AW_S3_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AW_S3_NMV 2
`define AXI_AW_S3_NMV_LOG2 1
`define AXI_AW_S3_NMV_P1_LOG2 2
`define AXI_W_S3_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_W_S3_NMV 2
`define AXI_W_S3_NMV_LOG2 1
`define AXI_W_S3_NMV_P1_LOG2 2
`define AXI_AR_S4_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AR_S4_NMV 1
`define AXI_AR_S4_NMV_LOG2 1
`define AXI_AR_S4_NMV_P1_LOG2 1
`define AXI_AW_S4_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AW_S4_NMV 1
`define AXI_AW_S4_NMV_LOG2 1
`define AXI_AW_S4_NMV_P1_LOG2 1
`define AXI_W_S4_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_W_S4_NMV 1
`define AXI_W_S4_NMV_LOG2 1
`define AXI_W_S4_NMV_P1_LOG2 1
`define AXI_AR_S5_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AR_S5_NMV 1
`define AXI_AR_S5_NMV_LOG2 1
`define AXI_AR_S5_NMV_P1_LOG2 1
`define AXI_AW_S5_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AW_S5_NMV 1
`define AXI_AW_S5_NMV_LOG2 1
`define AXI_AW_S5_NMV_P1_LOG2 1
`define AXI_W_S5_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_W_S5_NMV 1
`define AXI_W_S5_NMV_LOG2 1
`define AXI_W_S5_NMV_P1_LOG2 1
`define AXI_AR_S6_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AR_S6_NMV 1
`define AXI_AR_S6_NMV_LOG2 1
`define AXI_AR_S6_NMV_P1_LOG2 1
`define AXI_AW_S6_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AW_S6_NMV 1
`define AXI_AW_S6_NMV_LOG2 1
`define AXI_AW_S6_NMV_P1_LOG2 1
`define AXI_W_S6_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_W_S6_NMV 1
`define AXI_W_S6_NMV_LOG2 1
`define AXI_W_S6_NMV_P1_LOG2 1
`define AXI_AR_S7_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AR_S7_NMV 1
`define AXI_AR_S7_NMV_LOG2 1
`define AXI_AR_S7_NMV_P1_LOG2 1
`define AXI_AW_S7_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AW_S7_NMV 1
`define AXI_AW_S7_NMV_LOG2 1
`define AXI_AW_S7_NMV_P1_LOG2 1
`define AXI_W_S7_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_W_S7_NMV 1
`define AXI_W_S7_NMV_LOG2 1
`define AXI_W_S7_NMV_P1_LOG2 1
`define AXI_AR_S8_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AR_S8_NMV 1
`define AXI_AR_S8_NMV_LOG2 1
`define AXI_AR_S8_NMV_P1_LOG2 1
`define AXI_AW_S8_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AW_S8_NMV 1
`define AXI_AW_S8_NMV_LOG2 1
`define AXI_AW_S8_NMV_P1_LOG2 1
`define AXI_W_S8_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_W_S8_NMV 1
`define AXI_W_S8_NMV_LOG2 1
`define AXI_W_S8_NMV_P1_LOG2 1
`define AXI_AR_S9_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AR_S9_NMV 1
`define AXI_AR_S9_NMV_LOG2 1
`define AXI_AR_S9_NMV_P1_LOG2 1
`define AXI_AW_S9_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AW_S9_NMV 1
`define AXI_AW_S9_NMV_LOG2 1
`define AXI_AW_S9_NMV_P1_LOG2 1
`define AXI_W_S9_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_W_S9_NMV 1
`define AXI_W_S9_NMV_LOG2 1
`define AXI_W_S9_NMV_P1_LOG2 1
`define AXI_AR_S10_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AR_S10_NMV 1
`define AXI_AR_S10_NMV_LOG2 1
`define AXI_AR_S10_NMV_P1_LOG2 1
`define AXI_AW_S10_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AW_S10_NMV 1
`define AXI_AW_S10_NMV_LOG2 1
`define AXI_AW_S10_NMV_P1_LOG2 1
`define AXI_W_S10_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_W_S10_NMV 1
`define AXI_W_S10_NMV_LOG2 1
`define AXI_W_S10_NMV_P1_LOG2 1
`define AXI_AR_S11_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AR_S11_NMV 1
`define AXI_AR_S11_NMV_LOG2 1
`define AXI_AR_S11_NMV_P1_LOG2 1
`define AXI_AW_S11_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AW_S11_NMV 1
`define AXI_AW_S11_NMV_LOG2 1
`define AXI_AW_S11_NMV_P1_LOG2 1
`define AXI_W_S11_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_W_S11_NMV 1
`define AXI_W_S11_NMV_LOG2 1
`define AXI_W_S11_NMV_P1_LOG2 1
`define AXI_AR_S12_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AR_S12_NMV 1
`define AXI_AR_S12_NMV_LOG2 1
`define AXI_AR_S12_NMV_P1_LOG2 1
`define AXI_AW_S12_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AW_S12_NMV 1
`define AXI_AW_S12_NMV_LOG2 1
`define AXI_AW_S12_NMV_P1_LOG2 1
`define AXI_W_S12_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_W_S12_NMV 1
`define AXI_W_S12_NMV_LOG2 1
`define AXI_W_S12_NMV_P1_LOG2 1
`define AXI_AR_S13_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AR_S13_NMV 1
`define AXI_AR_S13_NMV_LOG2 1
`define AXI_AR_S13_NMV_P1_LOG2 1
`define AXI_AW_S13_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AW_S13_NMV 1
`define AXI_AW_S13_NMV_LOG2 1
`define AXI_AW_S13_NMV_P1_LOG2 1
`define AXI_W_S13_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_W_S13_NMV 1
`define AXI_W_S13_NMV_LOG2 1
`define AXI_W_S13_NMV_P1_LOG2 1
`define AXI_AR_S14_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AR_S14_NMV 1
`define AXI_AR_S14_NMV_LOG2 1
`define AXI_AR_S14_NMV_P1_LOG2 1
`define AXI_AW_S14_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AW_S14_NMV 1
`define AXI_AW_S14_NMV_LOG2 1
`define AXI_AW_S14_NMV_P1_LOG2 1
`define AXI_W_S14_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_W_S14_NMV 1
`define AXI_W_S14_NMV_LOG2 1
`define AXI_W_S14_NMV_P1_LOG2 1
`define AXI_AR_S15_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AR_S15_NMV 1
`define AXI_AR_S15_NMV_LOG2 1
`define AXI_AR_S15_NMV_P1_LOG2 1
`define AXI_AW_S15_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AW_S15_NMV 1
`define AXI_AW_S15_NMV_LOG2 1
`define AXI_AW_S15_NMV_P1_LOG2 1
`define AXI_W_S15_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_W_S15_NMV 1
`define AXI_W_S15_NMV_LOG2 1
`define AXI_W_S15_NMV_P1_LOG2 1
`define AXI_AR_S16_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AR_S16_NMV 1
`define AXI_AR_S16_NMV_LOG2 1
`define AXI_AR_S16_NMV_P1_LOG2 1
`define AXI_AW_S16_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_AW_S16_NMV 1
`define AXI_AW_S16_NMV_LOG2 1
`define AXI_AW_S16_NMV_P1_LOG2 1
`define AXI_W_S16_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_W_S16_NMV 1
`define AXI_W_S16_NMV_LOG2 1
`define AXI_W_S16_NMV_P1_LOG2 1
`define AXI_R_M1_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_R_M1_NSV 4
`define AXI_R_M1_NSV_LOG2 2
`define AXI_R_M1_NSV_P1_LOG2 3
`define AXI_B_M1_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_B_M1_NSV 4
`define AXI_B_M1_NSV_LOG2 2
`define AXI_B_M1_NSV_P1_LOG2 3
`define AXI_R_M2_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_R_M2_NSV 4
`define AXI_R_M2_NSV_LOG2 2
`define AXI_R_M2_NSV_P1_LOG2 3
`define AXI_B_M2_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_B_M2_NSV 4
`define AXI_B_M2_NSV_LOG2 2
`define AXI_B_M2_NSV_P1_LOG2 3
`define AXI_R_M3_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_R_M3_NSV 1
`define AXI_R_M3_NSV_LOG2 1
`define AXI_R_M3_NSV_P1_LOG2 1
`define AXI_B_M3_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_B_M3_NSV 1
`define AXI_B_M3_NSV_LOG2 1
`define AXI_B_M3_NSV_P1_LOG2 1
`define AXI_R_M4_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_R_M4_NSV 1
`define AXI_R_M4_NSV_LOG2 1
`define AXI_R_M4_NSV_P1_LOG2 1
`define AXI_B_M4_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_B_M4_NSV 1
`define AXI_B_M4_NSV_LOG2 1
`define AXI_B_M4_NSV_P1_LOG2 1
`define AXI_R_M5_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_R_M5_NSV 1
`define AXI_R_M5_NSV_LOG2 1
`define AXI_R_M5_NSV_P1_LOG2 1
`define AXI_B_M5_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_B_M5_NSV 1
`define AXI_B_M5_NSV_LOG2 1
`define AXI_B_M5_NSV_P1_LOG2 1
`define AXI_R_M6_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_R_M6_NSV 1
`define AXI_R_M6_NSV_LOG2 1
`define AXI_R_M6_NSV_P1_LOG2 1
`define AXI_B_M6_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_B_M6_NSV 1
`define AXI_B_M6_NSV_LOG2 1
`define AXI_B_M6_NSV_P1_LOG2 1
`define AXI_R_M7_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_R_M7_NSV 1
`define AXI_R_M7_NSV_LOG2 1
`define AXI_R_M7_NSV_P1_LOG2 1
`define AXI_B_M7_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_B_M7_NSV 1
`define AXI_B_M7_NSV_LOG2 1
`define AXI_B_M7_NSV_P1_LOG2 1
`define AXI_R_M8_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_R_M8_NSV 1
`define AXI_R_M8_NSV_LOG2 1
`define AXI_R_M8_NSV_P1_LOG2 1
`define AXI_B_M8_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_B_M8_NSV 1
`define AXI_B_M8_NSV_LOG2 1
`define AXI_B_M8_NSV_P1_LOG2 1
`define AXI_R_M9_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_R_M9_NSV 1
`define AXI_R_M9_NSV_LOG2 1
`define AXI_R_M9_NSV_P1_LOG2 1
`define AXI_B_M9_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_B_M9_NSV 1
`define AXI_B_M9_NSV_LOG2 1
`define AXI_B_M9_NSV_P1_LOG2 1
`define AXI_R_M10_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_R_M10_NSV 1
`define AXI_R_M10_NSV_LOG2 1
`define AXI_R_M10_NSV_P1_LOG2 1
`define AXI_B_M10_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_B_M10_NSV 1
`define AXI_B_M10_NSV_LOG2 1
`define AXI_B_M10_NSV_P1_LOG2 1
`define AXI_R_M11_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_R_M11_NSV 1
`define AXI_R_M11_NSV_LOG2 1
`define AXI_R_M11_NSV_P1_LOG2 1
`define AXI_B_M11_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_B_M11_NSV 1
`define AXI_B_M11_NSV_LOG2 1
`define AXI_B_M11_NSV_P1_LOG2 1
`define AXI_R_M12_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_R_M12_NSV 1
`define AXI_R_M12_NSV_LOG2 1
`define AXI_R_M12_NSV_P1_LOG2 1
`define AXI_B_M12_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_B_M12_NSV 1
`define AXI_B_M12_NSV_LOG2 1
`define AXI_B_M12_NSV_P1_LOG2 1
`define AXI_R_M13_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_R_M13_NSV 1
`define AXI_R_M13_NSV_LOG2 1
`define AXI_R_M13_NSV_P1_LOG2 1
`define AXI_B_M13_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_B_M13_NSV 1
`define AXI_B_M13_NSV_LOG2 1
`define AXI_B_M13_NSV_P1_LOG2 1
`define AXI_R_M14_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_R_M14_NSV 1
`define AXI_R_M14_NSV_LOG2 1
`define AXI_R_M14_NSV_P1_LOG2 1
`define AXI_B_M14_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_B_M14_NSV 1
`define AXI_B_M14_NSV_LOG2 1
`define AXI_B_M14_NSV_P1_LOG2 1
`define AXI_R_M15_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_R_M15_NSV 1
`define AXI_R_M15_NSV_LOG2 1
`define AXI_R_M15_NSV_P1_LOG2 1
`define AXI_B_M15_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_B_M15_NSV 1
`define AXI_B_M15_NSV_LOG2 1
`define AXI_B_M15_NSV_P1_LOG2 1
`define AXI_R_M16_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_R_M16_NSV 1
`define AXI_R_M16_NSV_LOG2 1
`define AXI_R_M16_NSV_P1_LOG2 1
`define AXI_B_M16_HAS_SHRD_DDCTD_LNK_VAL 0
`define AXI_B_M16_NSV 1
`define AXI_B_M16_NSV_LOG2 1
`define AXI_B_M16_NSV_P1_LOG2 1
`define AXI_M1_ON_AR_SHARED_VAL 0
`define AXI_M2_ON_AR_SHARED_VAL 0
`define AXI_M3_ON_AR_SHARED_VAL 0
`define AXI_M4_ON_AR_SHARED_VAL 0
`define AXI_M5_ON_AR_SHARED_VAL 0
`define AXI_M6_ON_AR_SHARED_VAL 0
`define AXI_M7_ON_AR_SHARED_VAL 0
`define AXI_M8_ON_AR_SHARED_VAL 0
`define AXI_M9_ON_AR_SHARED_VAL 0
`define AXI_M10_ON_AR_SHARED_VAL 0
`define AXI_M11_ON_AR_SHARED_VAL 0
`define AXI_M12_ON_AR_SHARED_VAL 0
`define AXI_M13_ON_AR_SHARED_VAL 0
`define AXI_M14_ON_AR_SHARED_VAL 0
`define AXI_M15_ON_AR_SHARED_VAL 0
`define AXI_M16_ON_AR_SHARED_VAL 0
`define AXI_S0_ON_AR_SHARED_VAL 0
`define AXI_S0_ON_AR_SHARED_ONLY_VAL 0
`define AXI_S1_ON_AR_SHARED_VAL 0
`define AXI_S1_ON_AR_SHARED_ONLY_VAL 0
`define AXI_S2_ON_AR_SHARED_VAL 0
`define AXI_S2_ON_AR_SHARED_ONLY_VAL 0
`define AXI_S3_ON_AR_SHARED_VAL 0
`define AXI_S3_ON_AR_SHARED_ONLY_VAL 0
`define AXI_S4_ON_AR_SHARED_VAL 0
`define AXI_S4_ON_AR_SHARED_ONLY
`define AXI_S4_ON_AR_SHARED_ONLY_VAL 1
`define AXI_S5_ON_AR_SHARED_VAL 0
`define AXI_S5_ON_AR_SHARED_ONLY
`define AXI_S5_ON_AR_SHARED_ONLY_VAL 1
`define AXI_S6_ON_AR_SHARED_VAL 0
`define AXI_S6_ON_AR_SHARED_ONLY
`define AXI_S6_ON_AR_SHARED_ONLY_VAL 1
`define AXI_S7_ON_AR_SHARED_VAL 0
`define AXI_S7_ON_AR_SHARED_ONLY
`define AXI_S7_ON_AR_SHARED_ONLY_VAL 1
`define AXI_S8_ON_AR_SHARED_VAL 0
`define AXI_S8_ON_AR_SHARED_ONLY
`define AXI_S8_ON_AR_SHARED_ONLY_VAL 1
`define AXI_S9_ON_AR_SHARED_VAL 0
`define AXI_S9_ON_AR_SHARED_ONLY
`define AXI_S9_ON_AR_SHARED_ONLY_VAL 1
`define AXI_S10_ON_AR_SHARED_VAL 0
`define AXI_S10_ON_AR_SHARED_ONLY
`define AXI_S10_ON_AR_SHARED_ONLY_VAL 1
`define AXI_S11_ON_AR_SHARED_VAL 0
`define AXI_S11_ON_AR_SHARED_ONLY
`define AXI_S11_ON_AR_SHARED_ONLY_VAL 1
`define AXI_S12_ON_AR_SHARED_VAL 0
`define AXI_S12_ON_AR_SHARED_ONLY
`define AXI_S12_ON_AR_SHARED_ONLY_VAL 1
`define AXI_S13_ON_AR_SHARED_VAL 0
`define AXI_S13_ON_AR_SHARED_ONLY
`define AXI_S13_ON_AR_SHARED_ONLY_VAL 1
`define AXI_S14_ON_AR_SHARED_VAL 0
`define AXI_S14_ON_AR_SHARED_ONLY
`define AXI_S14_ON_AR_SHARED_ONLY_VAL 1
`define AXI_S15_ON_AR_SHARED_VAL 0
`define AXI_S15_ON_AR_SHARED_ONLY
`define AXI_S15_ON_AR_SHARED_ONLY_VAL 1
`define AXI_S16_ON_AR_SHARED_VAL 0
`define AXI_S16_ON_AR_SHARED_ONLY
`define AXI_S16_ON_AR_SHARED_ONLY_VAL 1
`define AXI_M1_ON_AW_SHARED_VAL 0
`define AXI_M2_ON_AW_SHARED_VAL 0
`define AXI_M3_ON_AW_SHARED_VAL 0
`define AXI_M4_ON_AW_SHARED_VAL 0
`define AXI_M5_ON_AW_SHARED_VAL 0
`define AXI_M6_ON_AW_SHARED_VAL 0
`define AXI_M7_ON_AW_SHARED_VAL 0
`define AXI_M8_ON_AW_SHARED_VAL 0
`define AXI_M9_ON_AW_SHARED_VAL 0
`define AXI_M10_ON_AW_SHARED_VAL 0
`define AXI_M11_ON_AW_SHARED_VAL 0
`define AXI_M12_ON_AW_SHARED_VAL 0
`define AXI_M13_ON_AW_SHARED_VAL 0
`define AXI_M14_ON_AW_SHARED_VAL 0
`define AXI_M15_ON_AW_SHARED_VAL 0
`define AXI_M16_ON_AW_SHARED_VAL 0
`define AXI_S0_ON_AW_SHARED_VAL 0
`define AXI_S0_ON_AW_SHARED_ONLY_VAL 0
`define AXI_S1_ON_AW_SHARED_VAL 0
`define AXI_S1_ON_AW_SHARED_ONLY_VAL 0
`define AXI_S2_ON_AW_SHARED_VAL 0
`define AXI_S2_ON_AW_SHARED_ONLY_VAL 0
`define AXI_S3_ON_AW_SHARED_VAL 0
`define AXI_S3_ON_AW_SHARED_ONLY_VAL 0
`define AXI_S4_ON_AW_SHARED_VAL 0
`define AXI_S4_ON_AW_SHARED_ONLY
`define AXI_S4_ON_AW_SHARED_ONLY_VAL 1
`define AXI_S5_ON_AW_SHARED_VAL 0
`define AXI_S5_ON_AW_SHARED_ONLY
`define AXI_S5_ON_AW_SHARED_ONLY_VAL 1
`define AXI_S6_ON_AW_SHARED_VAL 0
`define AXI_S6_ON_AW_SHARED_ONLY
`define AXI_S6_ON_AW_SHARED_ONLY_VAL 1
`define AXI_S7_ON_AW_SHARED_VAL 0
`define AXI_S7_ON_AW_SHARED_ONLY
`define AXI_S7_ON_AW_SHARED_ONLY_VAL 1
`define AXI_S8_ON_AW_SHARED_VAL 0
`define AXI_S8_ON_AW_SHARED_ONLY
`define AXI_S8_ON_AW_SHARED_ONLY_VAL 1
`define AXI_S9_ON_AW_SHARED_VAL 0
`define AXI_S9_ON_AW_SHARED_ONLY
`define AXI_S9_ON_AW_SHARED_ONLY_VAL 1
`define AXI_S10_ON_AW_SHARED_VAL 0
`define AXI_S10_ON_AW_SHARED_ONLY
`define AXI_S10_ON_AW_SHARED_ONLY_VAL 1
`define AXI_S11_ON_AW_SHARED_VAL 0
`define AXI_S11_ON_AW_SHARED_ONLY
`define AXI_S11_ON_AW_SHARED_ONLY_VAL 1
`define AXI_S12_ON_AW_SHARED_VAL 0
`define AXI_S12_ON_AW_SHARED_ONLY
`define AXI_S12_ON_AW_SHARED_ONLY_VAL 1
`define AXI_S13_ON_AW_SHARED_VAL 0
`define AXI_S13_ON_AW_SHARED_ONLY
`define AXI_S13_ON_AW_SHARED_ONLY_VAL 1
`define AXI_S14_ON_AW_SHARED_VAL 0
`define AXI_S14_ON_AW_SHARED_ONLY
`define AXI_S14_ON_AW_SHARED_ONLY_VAL 1
`define AXI_S15_ON_AW_SHARED_VAL 0
`define AXI_S15_ON_AW_SHARED_ONLY
`define AXI_S15_ON_AW_SHARED_ONLY_VAL 1
`define AXI_S16_ON_AW_SHARED_VAL 0
`define AXI_S16_ON_AW_SHARED_ONLY
`define AXI_S16_ON_AW_SHARED_ONLY_VAL 1
`define AXI_M1_ON_W_SHARED_VAL 0
`define AXI_M2_ON_W_SHARED_VAL 0
`define AXI_M3_ON_W_SHARED_VAL 0
`define AXI_M4_ON_W_SHARED_VAL 0
`define AXI_M5_ON_W_SHARED_VAL 0
`define AXI_M6_ON_W_SHARED_VAL 0
`define AXI_M7_ON_W_SHARED_VAL 0
`define AXI_M8_ON_W_SHARED_VAL 0
`define AXI_M9_ON_W_SHARED_VAL 0
`define AXI_M10_ON_W_SHARED_VAL 0
`define AXI_M11_ON_W_SHARED_VAL 0
`define AXI_M12_ON_W_SHARED_VAL 0
`define AXI_M13_ON_W_SHARED_VAL 0
`define AXI_M14_ON_W_SHARED_VAL 0
`define AXI_M15_ON_W_SHARED_VAL 0
`define AXI_M16_ON_W_SHARED_VAL 0
`define AXI_S0_ON_W_SHARED_VAL 0
`define AXI_S0_ON_W_SHARED_ONLY_VAL 0
`define AXI_S1_ON_W_SHARED_VAL 0
`define AXI_S1_ON_W_SHARED_ONLY_VAL 0
`define AXI_S2_ON_W_SHARED_VAL 0
`define AXI_S2_ON_W_SHARED_ONLY_VAL 0
`define AXI_S3_ON_W_SHARED_VAL 0
`define AXI_S3_ON_W_SHARED_ONLY_VAL 0
`define AXI_S4_ON_W_SHARED_VAL 0
`define AXI_S4_ON_W_SHARED_ONLY
`define AXI_S4_ON_W_SHARED_ONLY_VAL 1
`define AXI_S5_ON_W_SHARED_VAL 0
`define AXI_S5_ON_W_SHARED_ONLY
`define AXI_S5_ON_W_SHARED_ONLY_VAL 1
`define AXI_S6_ON_W_SHARED_VAL 0
`define AXI_S6_ON_W_SHARED_ONLY
`define AXI_S6_ON_W_SHARED_ONLY_VAL 1
`define AXI_S7_ON_W_SHARED_VAL 0
`define AXI_S7_ON_W_SHARED_ONLY
`define AXI_S7_ON_W_SHARED_ONLY_VAL 1
`define AXI_S8_ON_W_SHARED_VAL 0
`define AXI_S8_ON_W_SHARED_ONLY
`define AXI_S8_ON_W_SHARED_ONLY_VAL 1
`define AXI_S9_ON_W_SHARED_VAL 0
`define AXI_S9_ON_W_SHARED_ONLY
`define AXI_S9_ON_W_SHARED_ONLY_VAL 1
`define AXI_S10_ON_W_SHARED_VAL 0
`define AXI_S10_ON_W_SHARED_ONLY
`define AXI_S10_ON_W_SHARED_ONLY_VAL 1
`define AXI_S11_ON_W_SHARED_VAL 0
`define AXI_S11_ON_W_SHARED_ONLY
`define AXI_S11_ON_W_SHARED_ONLY_VAL 1
`define AXI_S12_ON_W_SHARED_VAL 0
`define AXI_S12_ON_W_SHARED_ONLY
`define AXI_S12_ON_W_SHARED_ONLY_VAL 1
`define AXI_S13_ON_W_SHARED_VAL 0
`define AXI_S13_ON_W_SHARED_ONLY
`define AXI_S13_ON_W_SHARED_ONLY_VAL 1
`define AXI_S14_ON_W_SHARED_VAL 0
`define AXI_S14_ON_W_SHARED_ONLY
`define AXI_S14_ON_W_SHARED_ONLY_VAL 1
`define AXI_S15_ON_W_SHARED_VAL 0
`define AXI_S15_ON_W_SHARED_ONLY
`define AXI_S15_ON_W_SHARED_ONLY_VAL 1
`define AXI_S16_ON_W_SHARED_VAL 0
`define AXI_S16_ON_W_SHARED_ONLY
`define AXI_S16_ON_W_SHARED_ONLY_VAL 1
`define AXI_S0_ON_R_SHARED_VAL 0
`define AXI_S1_ON_R_SHARED_VAL 0
`define AXI_S2_ON_R_SHARED_VAL 0
`define AXI_S3_ON_R_SHARED_VAL 0
`define AXI_S4_ON_R_SHARED_VAL 0
`define AXI_S5_ON_R_SHARED_VAL 0
`define AXI_S6_ON_R_SHARED_VAL 0
`define AXI_S7_ON_R_SHARED_VAL 0
`define AXI_S8_ON_R_SHARED_VAL 0
`define AXI_S9_ON_R_SHARED_VAL 0
`define AXI_S10_ON_R_SHARED_VAL 0
`define AXI_S11_ON_R_SHARED_VAL 0
`define AXI_S12_ON_R_SHARED_VAL 0
`define AXI_S13_ON_R_SHARED_VAL 0
`define AXI_S14_ON_R_SHARED_VAL 0
`define AXI_S15_ON_R_SHARED_VAL 0
`define AXI_S16_ON_R_SHARED_VAL 0
`define AXI_M1_ON_R_SHARED_VAL 0
`define AXI_M1_ON_R_SHARED_ONLY_VAL 0
`define AXI_M2_ON_R_SHARED_VAL 0
`define AXI_M2_ON_R_SHARED_ONLY_VAL 0
`define AXI_M3_ON_R_SHARED_VAL 0
`define AXI_M3_ON_R_SHARED_ONLY
`define AXI_M3_ON_R_SHARED_ONLY_VAL 1
`define AXI_M4_ON_R_SHARED_VAL 0
`define AXI_M4_ON_R_SHARED_ONLY
`define AXI_M4_ON_R_SHARED_ONLY_VAL 1
`define AXI_M5_ON_R_SHARED_VAL 0
`define AXI_M5_ON_R_SHARED_ONLY
`define AXI_M5_ON_R_SHARED_ONLY_VAL 1
`define AXI_M6_ON_R_SHARED_VAL 0
`define AXI_M6_ON_R_SHARED_ONLY
`define AXI_M6_ON_R_SHARED_ONLY_VAL 1
`define AXI_M7_ON_R_SHARED_VAL 0
`define AXI_M7_ON_R_SHARED_ONLY
`define AXI_M7_ON_R_SHARED_ONLY_VAL 1
`define AXI_M8_ON_R_SHARED_VAL 0
`define AXI_M8_ON_R_SHARED_ONLY
`define AXI_M8_ON_R_SHARED_ONLY_VAL 1
`define AXI_M9_ON_R_SHARED_VAL 0
`define AXI_M9_ON_R_SHARED_ONLY
`define AXI_M9_ON_R_SHARED_ONLY_VAL 1
`define AXI_M10_ON_R_SHARED_VAL 0
`define AXI_M10_ON_R_SHARED_ONLY
`define AXI_M10_ON_R_SHARED_ONLY_VAL 1
`define AXI_M11_ON_R_SHARED_VAL 0
`define AXI_M11_ON_R_SHARED_ONLY
`define AXI_M11_ON_R_SHARED_ONLY_VAL 1
`define AXI_M12_ON_R_SHARED_VAL 0
`define AXI_M12_ON_R_SHARED_ONLY
`define AXI_M12_ON_R_SHARED_ONLY_VAL 1
`define AXI_M13_ON_R_SHARED_VAL 0
`define AXI_M13_ON_R_SHARED_ONLY
`define AXI_M13_ON_R_SHARED_ONLY_VAL 1
`define AXI_M14_ON_R_SHARED_VAL 0
`define AXI_M14_ON_R_SHARED_ONLY
`define AXI_M14_ON_R_SHARED_ONLY_VAL 1
`define AXI_M15_ON_R_SHARED_VAL 0
`define AXI_M15_ON_R_SHARED_ONLY
`define AXI_M15_ON_R_SHARED_ONLY_VAL 1
`define AXI_M16_ON_R_SHARED_VAL 0
`define AXI_M16_ON_R_SHARED_ONLY
`define AXI_M16_ON_R_SHARED_ONLY_VAL 1
`define AXI_S0_ON_B_SHARED_VAL 0
`define AXI_S1_ON_B_SHARED_VAL 0
`define AXI_S2_ON_B_SHARED_VAL 0
`define AXI_S3_ON_B_SHARED_VAL 0
`define AXI_S4_ON_B_SHARED_VAL 0
`define AXI_S5_ON_B_SHARED_VAL 0
`define AXI_S6_ON_B_SHARED_VAL 0
`define AXI_S7_ON_B_SHARED_VAL 0
`define AXI_S8_ON_B_SHARED_VAL 0
`define AXI_S9_ON_B_SHARED_VAL 0
`define AXI_S10_ON_B_SHARED_VAL 0
`define AXI_S11_ON_B_SHARED_VAL 0
`define AXI_S12_ON_B_SHARED_VAL 0
`define AXI_S13_ON_B_SHARED_VAL 0
`define AXI_S14_ON_B_SHARED_VAL 0
`define AXI_S15_ON_B_SHARED_VAL 0
`define AXI_S16_ON_B_SHARED_VAL 0
`define AXI_M1_ON_B_SHARED_VAL 0
`define AXI_M1_ON_B_SHARED_ONLY_VAL 0
`define AXI_M2_ON_B_SHARED_VAL 0
`define AXI_M2_ON_B_SHARED_ONLY_VAL 0
`define AXI_M3_ON_B_SHARED_VAL 0
`define AXI_M3_ON_B_SHARED_ONLY
`define AXI_M3_ON_B_SHARED_ONLY_VAL 1
`define AXI_M4_ON_B_SHARED_VAL 0
`define AXI_M4_ON_B_SHARED_ONLY
`define AXI_M4_ON_B_SHARED_ONLY_VAL 1
`define AXI_M5_ON_B_SHARED_VAL 0
`define AXI_M5_ON_B_SHARED_ONLY
`define AXI_M5_ON_B_SHARED_ONLY_VAL 1
`define AXI_M6_ON_B_SHARED_VAL 0
`define AXI_M6_ON_B_SHARED_ONLY
`define AXI_M6_ON_B_SHARED_ONLY_VAL 1
`define AXI_M7_ON_B_SHARED_VAL 0
`define AXI_M7_ON_B_SHARED_ONLY
`define AXI_M7_ON_B_SHARED_ONLY_VAL 1
`define AXI_M8_ON_B_SHARED_VAL 0
`define AXI_M8_ON_B_SHARED_ONLY
`define AXI_M8_ON_B_SHARED_ONLY_VAL 1
`define AXI_M9_ON_B_SHARED_VAL 0
`define AXI_M9_ON_B_SHARED_ONLY
`define AXI_M9_ON_B_SHARED_ONLY_VAL 1
`define AXI_M10_ON_B_SHARED_VAL 0
`define AXI_M10_ON_B_SHARED_ONLY
`define AXI_M10_ON_B_SHARED_ONLY_VAL 1
`define AXI_M11_ON_B_SHARED_VAL 0
`define AXI_M11_ON_B_SHARED_ONLY
`define AXI_M11_ON_B_SHARED_ONLY_VAL 1
`define AXI_M12_ON_B_SHARED_VAL 0
`define AXI_M12_ON_B_SHARED_ONLY
`define AXI_M12_ON_B_SHARED_ONLY_VAL 1
`define AXI_M13_ON_B_SHARED_VAL 0
`define AXI_M13_ON_B_SHARED_ONLY
`define AXI_M13_ON_B_SHARED_ONLY_VAL 1
`define AXI_M14_ON_B_SHARED_VAL 0
`define AXI_M14_ON_B_SHARED_ONLY
`define AXI_M14_ON_B_SHARED_ONLY_VAL 1
`define AXI_M15_ON_B_SHARED_VAL 0
`define AXI_M15_ON_B_SHARED_ONLY
`define AXI_M15_ON_B_SHARED_ONLY_VAL 1
`define AXI_M16_ON_B_SHARED_VAL 0
`define AXI_M16_ON_B_SHARED_ONLY
`define AXI_M16_ON_B_SHARED_ONLY_VAL 1
`define AXI_AW_SHARED_PL 0
`define AXI_AR_SHARED_PL 0
`define AXI_W_SHARED_PL 0
`define AXI_R_SHARED_PL 0
`define AXI_B_SHARED_PL 0
`define AXI_MCA_HLD_PRIOR 0
`define AXI_AR_MCA_NC_S0 1
`define AXI_AR_MCA_EN_S0 (`AXI_AR_MCA_NC_S0 > 1)
`define AXI_AR_MCA_NC_W_S0 1
`define AXI_AW_MCA_NC_S0 1
`define AXI_AW_MCA_EN_S0 (`AXI_AW_MCA_NC_S0 > 1)
`define AXI_AW_MCA_NC_W_S0 1
`define AXI_W_MCA_NC_S0 1
`define AXI_W_MCA_EN_S0 (`AXI_W_MCA_NC_S0 > 1)
`define AXI_W_MCA_NC_W_S0 1
`define AXI_AR_MCA_NC_S1 1
`define AXI_AR_MCA_EN_S1 (`AXI_AR_MCA_NC_S1 > 1)
`define AXI_AR_MCA_NC_W_S1 1
`define AXI_AW_MCA_NC_S1 1
`define AXI_AW_MCA_EN_S1 (`AXI_AW_MCA_NC_S1 > 1)
`define AXI_AW_MCA_NC_W_S1 1
`define AXI_W_MCA_NC_S1 1
`define AXI_W_MCA_EN_S1 (`AXI_W_MCA_NC_S1 > 1)
`define AXI_W_MCA_NC_W_S1 1
`define AXI_AR_MCA_NC_S2 1
`define AXI_AR_MCA_EN_S2 (`AXI_AR_MCA_NC_S2 > 1)
`define AXI_AR_MCA_NC_W_S2 1
`define AXI_AW_MCA_NC_S2 1
`define AXI_AW_MCA_EN_S2 (`AXI_AW_MCA_NC_S2 > 1)
`define AXI_AW_MCA_NC_W_S2 1
`define AXI_W_MCA_NC_S2 1
`define AXI_W_MCA_EN_S2 (`AXI_W_MCA_NC_S2 > 1)
`define AXI_W_MCA_NC_W_S2 1
`define AXI_AR_MCA_NC_S3 1
`define AXI_AR_MCA_EN_S3 (`AXI_AR_MCA_NC_S3 > 1)
`define AXI_AR_MCA_NC_W_S3 1
`define AXI_AW_MCA_NC_S3 1
`define AXI_AW_MCA_EN_S3 (`AXI_AW_MCA_NC_S3 > 1)
`define AXI_AW_MCA_NC_W_S3 1
`define AXI_W_MCA_NC_S3 1
`define AXI_W_MCA_EN_S3 (`AXI_W_MCA_NC_S3 > 1)
`define AXI_W_MCA_NC_W_S3 1
`define AXI_AR_MCA_NC_S4 1
`define AXI_AR_MCA_EN_S4 (`AXI_AR_MCA_NC_S4 > 1)
`define AXI_AR_MCA_NC_W_S4 1
`define AXI_AW_MCA_NC_S4 1
`define AXI_AW_MCA_EN_S4 (`AXI_AW_MCA_NC_S4 > 1)
`define AXI_AW_MCA_NC_W_S4 1
`define AXI_W_MCA_NC_S4 1
`define AXI_W_MCA_EN_S4 (`AXI_W_MCA_NC_S4 > 1)
`define AXI_W_MCA_NC_W_S4 1
`define AXI_AR_MCA_NC_S5 1
`define AXI_AR_MCA_EN_S5 (`AXI_AR_MCA_NC_S5 > 1)
`define AXI_AR_MCA_NC_W_S5 1
`define AXI_AW_MCA_NC_S5 1
`define AXI_AW_MCA_EN_S5 (`AXI_AW_MCA_NC_S5 > 1)
`define AXI_AW_MCA_NC_W_S5 1
`define AXI_W_MCA_NC_S5 1
`define AXI_W_MCA_EN_S5 (`AXI_W_MCA_NC_S5 > 1)
`define AXI_W_MCA_NC_W_S5 1
`define AXI_AR_MCA_NC_S6 1
`define AXI_AR_MCA_EN_S6 (`AXI_AR_MCA_NC_S6 > 1)
`define AXI_AR_MCA_NC_W_S6 1
`define AXI_AW_MCA_NC_S6 1
`define AXI_AW_MCA_EN_S6 (`AXI_AW_MCA_NC_S6 > 1)
`define AXI_AW_MCA_NC_W_S6 1
`define AXI_W_MCA_NC_S6 1
`define AXI_W_MCA_EN_S6 (`AXI_W_MCA_NC_S6 > 1)
`define AXI_W_MCA_NC_W_S6 1
`define AXI_AR_MCA_NC_S7 1
`define AXI_AR_MCA_EN_S7 (`AXI_AR_MCA_NC_S7 > 1)
`define AXI_AR_MCA_NC_W_S7 1
`define AXI_AW_MCA_NC_S7 1
`define AXI_AW_MCA_EN_S7 (`AXI_AW_MCA_NC_S7 > 1)
`define AXI_AW_MCA_NC_W_S7 1
`define AXI_W_MCA_NC_S7 1
`define AXI_W_MCA_EN_S7 (`AXI_W_MCA_NC_S7 > 1)
`define AXI_W_MCA_NC_W_S7 1
`define AXI_AR_MCA_NC_S8 1
`define AXI_AR_MCA_EN_S8 (`AXI_AR_MCA_NC_S8 > 1)
`define AXI_AR_MCA_NC_W_S8 1
`define AXI_AW_MCA_NC_S8 1
`define AXI_AW_MCA_EN_S8 (`AXI_AW_MCA_NC_S8 > 1)
`define AXI_AW_MCA_NC_W_S8 1
`define AXI_W_MCA_NC_S8 1
`define AXI_W_MCA_EN_S8 (`AXI_W_MCA_NC_S8 > 1)
`define AXI_W_MCA_NC_W_S8 1
`define AXI_AR_MCA_NC_S9 1
`define AXI_AR_MCA_EN_S9 (`AXI_AR_MCA_NC_S9 > 1)
`define AXI_AR_MCA_NC_W_S9 1
`define AXI_AW_MCA_NC_S9 1
`define AXI_AW_MCA_EN_S9 (`AXI_AW_MCA_NC_S9 > 1)
`define AXI_AW_MCA_NC_W_S9 1
`define AXI_W_MCA_NC_S9 1
`define AXI_W_MCA_EN_S9 (`AXI_W_MCA_NC_S9 > 1)
`define AXI_W_MCA_NC_W_S9 1
`define AXI_AR_MCA_NC_S10 1
`define AXI_AR_MCA_EN_S10 (`AXI_AR_MCA_NC_S10 > 1)
`define AXI_AR_MCA_NC_W_S10 1
`define AXI_AW_MCA_NC_S10 1
`define AXI_AW_MCA_EN_S10 (`AXI_AW_MCA_NC_S10 > 1)
`define AXI_AW_MCA_NC_W_S10 1
`define AXI_W_MCA_NC_S10 1
`define AXI_W_MCA_EN_S10 (`AXI_W_MCA_NC_S10 > 1)
`define AXI_W_MCA_NC_W_S10 1
`define AXI_AR_MCA_NC_S11 1
`define AXI_AR_MCA_EN_S11 (`AXI_AR_MCA_NC_S11 > 1)
`define AXI_AR_MCA_NC_W_S11 1
`define AXI_AW_MCA_NC_S11 1
`define AXI_AW_MCA_EN_S11 (`AXI_AW_MCA_NC_S11 > 1)
`define AXI_AW_MCA_NC_W_S11 1
`define AXI_W_MCA_NC_S11 1
`define AXI_W_MCA_EN_S11 (`AXI_W_MCA_NC_S11 > 1)
`define AXI_W_MCA_NC_W_S11 1
`define AXI_AR_MCA_NC_S12 1
`define AXI_AR_MCA_EN_S12 (`AXI_AR_MCA_NC_S12 > 1)
`define AXI_AR_MCA_NC_W_S12 1
`define AXI_AW_MCA_NC_S12 1
`define AXI_AW_MCA_EN_S12 (`AXI_AW_MCA_NC_S12 > 1)
`define AXI_AW_MCA_NC_W_S12 1
`define AXI_W_MCA_NC_S12 1
`define AXI_W_MCA_EN_S12 (`AXI_W_MCA_NC_S12 > 1)
`define AXI_W_MCA_NC_W_S12 1
`define AXI_AR_MCA_NC_S13 1
`define AXI_AR_MCA_EN_S13 (`AXI_AR_MCA_NC_S13 > 1)
`define AXI_AR_MCA_NC_W_S13 1
`define AXI_AW_MCA_NC_S13 1
`define AXI_AW_MCA_EN_S13 (`AXI_AW_MCA_NC_S13 > 1)
`define AXI_AW_MCA_NC_W_S13 1
`define AXI_W_MCA_NC_S13 1
`define AXI_W_MCA_EN_S13 (`AXI_W_MCA_NC_S13 > 1)
`define AXI_W_MCA_NC_W_S13 1
`define AXI_AR_MCA_NC_S14 1
`define AXI_AR_MCA_EN_S14 (`AXI_AR_MCA_NC_S14 > 1)
`define AXI_AR_MCA_NC_W_S14 1
`define AXI_AW_MCA_NC_S14 1
`define AXI_AW_MCA_EN_S14 (`AXI_AW_MCA_NC_S14 > 1)
`define AXI_AW_MCA_NC_W_S14 1
`define AXI_W_MCA_NC_S14 1
`define AXI_W_MCA_EN_S14 (`AXI_W_MCA_NC_S14 > 1)
`define AXI_W_MCA_NC_W_S14 1
`define AXI_AR_MCA_NC_S15 1
`define AXI_AR_MCA_EN_S15 (`AXI_AR_MCA_NC_S15 > 1)
`define AXI_AR_MCA_NC_W_S15 1
`define AXI_AW_MCA_NC_S15 1
`define AXI_AW_MCA_EN_S15 (`AXI_AW_MCA_NC_S15 > 1)
`define AXI_AW_MCA_NC_W_S15 1
`define AXI_W_MCA_NC_S15 1
`define AXI_W_MCA_EN_S15 (`AXI_W_MCA_NC_S15 > 1)
`define AXI_W_MCA_NC_W_S15 1
`define AXI_AR_MCA_NC_S16 1
`define AXI_AR_MCA_EN_S16 (`AXI_AR_MCA_NC_S16 > 1)
`define AXI_AR_MCA_NC_W_S16 1
`define AXI_AW_MCA_NC_S16 1
`define AXI_AW_MCA_EN_S16 (`AXI_AW_MCA_NC_S16 > 1)
`define AXI_AW_MCA_NC_W_S16 1
`define AXI_W_MCA_NC_S16 1
`define AXI_W_MCA_EN_S16 (`AXI_W_MCA_NC_S16 > 1)
`define AXI_W_MCA_NC_W_S16 1
`define AXI_R_MCA_NC_M1 1
`define AXI_R_MCA_EN_M1 (`AXI_R_MCA_NC_M1 > 1)
`define AXI_R_MCA_NC_W_M1 1
`define AXI_B_MCA_NC_M1 1
`define AXI_B_MCA_EN_M1 (`AXI_B_MCA_NC_M1 > 1)
`define AXI_B_MCA_NC_W_M1 1
`define AXI_R_MCA_NC_M2 1
`define AXI_R_MCA_EN_M2 (`AXI_R_MCA_NC_M2 > 1)
`define AXI_R_MCA_NC_W_M2 1
`define AXI_B_MCA_NC_M2 1
`define AXI_B_MCA_EN_M2 (`AXI_B_MCA_NC_M2 > 1)
`define AXI_B_MCA_NC_W_M2 1
`define AXI_R_MCA_NC_M3 1
`define AXI_R_MCA_EN_M3 (`AXI_R_MCA_NC_M3 > 1)
`define AXI_R_MCA_NC_W_M3 1
`define AXI_B_MCA_NC_M3 1
`define AXI_B_MCA_EN_M3 (`AXI_B_MCA_NC_M3 > 1)
`define AXI_B_MCA_NC_W_M3 1
`define AXI_R_MCA_NC_M4 1
`define AXI_R_MCA_EN_M4 (`AXI_R_MCA_NC_M4 > 1)
`define AXI_R_MCA_NC_W_M4 1
`define AXI_B_MCA_NC_M4 1
`define AXI_B_MCA_EN_M4 (`AXI_B_MCA_NC_M4 > 1)
`define AXI_B_MCA_NC_W_M4 1
`define AXI_R_MCA_NC_M5 1
`define AXI_R_MCA_EN_M5 (`AXI_R_MCA_NC_M5 > 1)
`define AXI_R_MCA_NC_W_M5 1
`define AXI_B_MCA_NC_M5 1
`define AXI_B_MCA_EN_M5 (`AXI_B_MCA_NC_M5 > 1)
`define AXI_B_MCA_NC_W_M5 1
`define AXI_R_MCA_NC_M6 1
`define AXI_R_MCA_EN_M6 (`AXI_R_MCA_NC_M6 > 1)
`define AXI_R_MCA_NC_W_M6 1
`define AXI_B_MCA_NC_M6 1
`define AXI_B_MCA_EN_M6 (`AXI_B_MCA_NC_M6 > 1)
`define AXI_B_MCA_NC_W_M6 1
`define AXI_R_MCA_NC_M7 1
`define AXI_R_MCA_EN_M7 (`AXI_R_MCA_NC_M7 > 1)
`define AXI_R_MCA_NC_W_M7 1
`define AXI_B_MCA_NC_M7 1
`define AXI_B_MCA_EN_M7 (`AXI_B_MCA_NC_M7 > 1)
`define AXI_B_MCA_NC_W_M7 1
`define AXI_R_MCA_NC_M8 1
`define AXI_R_MCA_EN_M8 (`AXI_R_MCA_NC_M8 > 1)
`define AXI_R_MCA_NC_W_M8 1
`define AXI_B_MCA_NC_M8 1
`define AXI_B_MCA_EN_M8 (`AXI_B_MCA_NC_M8 > 1)
`define AXI_B_MCA_NC_W_M8 1
`define AXI_R_MCA_NC_M9 1
`define AXI_R_MCA_EN_M9 (`AXI_R_MCA_NC_M9 > 1)
`define AXI_R_MCA_NC_W_M9 1
`define AXI_B_MCA_NC_M9 1
`define AXI_B_MCA_EN_M9 (`AXI_B_MCA_NC_M9 > 1)
`define AXI_B_MCA_NC_W_M9 1
`define AXI_R_MCA_NC_M10 1
`define AXI_R_MCA_EN_M10 (`AXI_R_MCA_NC_M10 > 1)
`define AXI_R_MCA_NC_W_M10 1
`define AXI_B_MCA_NC_M10 1
`define AXI_B_MCA_EN_M10 (`AXI_B_MCA_NC_M10 > 1)
`define AXI_B_MCA_NC_W_M10 1
`define AXI_R_MCA_NC_M11 1
`define AXI_R_MCA_EN_M11 (`AXI_R_MCA_NC_M11 > 1)
`define AXI_R_MCA_NC_W_M11 1
`define AXI_B_MCA_NC_M11 1
`define AXI_B_MCA_EN_M11 (`AXI_B_MCA_NC_M11 > 1)
`define AXI_B_MCA_NC_W_M11 1
`define AXI_R_MCA_NC_M12 1
`define AXI_R_MCA_EN_M12 (`AXI_R_MCA_NC_M12 > 1)
`define AXI_R_MCA_NC_W_M12 1
`define AXI_B_MCA_NC_M12 1
`define AXI_B_MCA_EN_M12 (`AXI_B_MCA_NC_M12 > 1)
`define AXI_B_MCA_NC_W_M12 1
`define AXI_R_MCA_NC_M13 1
`define AXI_R_MCA_EN_M13 (`AXI_R_MCA_NC_M13 > 1)
`define AXI_R_MCA_NC_W_M13 1
`define AXI_B_MCA_NC_M13 1
`define AXI_B_MCA_EN_M13 (`AXI_B_MCA_NC_M13 > 1)
`define AXI_B_MCA_NC_W_M13 1
`define AXI_R_MCA_NC_M14 1
`define AXI_R_MCA_EN_M14 (`AXI_R_MCA_NC_M14 > 1)
`define AXI_R_MCA_NC_W_M14 1
`define AXI_B_MCA_NC_M14 1
`define AXI_B_MCA_EN_M14 (`AXI_B_MCA_NC_M14 > 1)
`define AXI_B_MCA_NC_W_M14 1
`define AXI_R_MCA_NC_M15 1
`define AXI_R_MCA_EN_M15 (`AXI_R_MCA_NC_M15 > 1)
`define AXI_R_MCA_NC_W_M15 1
`define AXI_B_MCA_NC_M15 1
`define AXI_B_MCA_EN_M15 (`AXI_B_MCA_NC_M15 > 1)
`define AXI_B_MCA_NC_W_M15 1
`define AXI_R_MCA_NC_M16 1
`define AXI_R_MCA_EN_M16 (`AXI_R_MCA_NC_M16 > 1)
`define AXI_R_MCA_NC_W_M16 1
`define AXI_B_MCA_NC_M16 1
`define AXI_B_MCA_EN_M16 (`AXI_B_MCA_NC_M16 > 1)
`define AXI_B_MCA_NC_W_M16 1
`define AXI_AR_SHARED_MCA_NC 1
`define AXI_AR_SHARED_MCA_EN (`AXI_AR_SHARED_MCA_NC > 1)
`define AXI_AR_SHARED_MCA_NC_W 1
`define AXI_AW_SHARED_MCA_NC 1
`define AXI_AW_SHARED_MCA_EN (`AXI_AW_SHARED_MCA_NC > 1)
`define AXI_AW_SHARED_MCA_NC_W 1
`define AXI_W_SHARED_MCA_NC 1
`define AXI_W_SHARED_MCA_EN (`AXI_W_SHARED_MCA_NC > 1)
`define AXI_W_SHARED_MCA_NC_W 1
`define AXI_R_SHARED_MCA_NC 1
`define AXI_R_SHARED_MCA_EN (`AXI_R_SHARED_MCA_NC > 1) 
`define AXI_R_SHARED_MCA_NC_W 1
`define AXI_B_SHARED_MCA_NC 1
`define AXI_B_SHARED_MCA_EN (`AXI_B_SHARED_MCA_NC > 1) 
`define AXI_B_SHARED_MCA_NC_W 1
`define AXI_MAX_RCA_ID_M1 4
`define AXI_LOG2_MAX_RCA_ID_P1_M1 3
`define AXI_MAX_WCA_ID_M1 4
`define AXI_LOG2_MAX_WCA_ID_P1_M1 3
`define AXI_MAX_URIDA_M1 5
`define AXI_LOG2_MAX_URIDA_M1 3
`define AXI_MAX_UWIDA_M1 5
`define AXI_LOG2_MAX_UWIDA_M1 3
`define AXI_RI_LIMIT_M1 0
`define AXI_MAX_RCA_ID_M2 4
`define AXI_LOG2_MAX_RCA_ID_P1_M2 3
`define AXI_MAX_WCA_ID_M2 4
`define AXI_LOG2_MAX_WCA_ID_P1_M2 3
`define AXI_MAX_URIDA_M2 5
`define AXI_LOG2_MAX_URIDA_M2 3
`define AXI_MAX_UWIDA_M2 5
`define AXI_LOG2_MAX_UWIDA_M2 3
`define AXI_RI_LIMIT_M2 0
`define AXI_MAX_RCA_ID_M3 4
`define AXI_LOG2_MAX_RCA_ID_P1_M3 3
`define AXI_MAX_WCA_ID_M3 4
`define AXI_LOG2_MAX_WCA_ID_P1_M3 3
`define AXI_MAX_URIDA_M3 5
`define AXI_LOG2_MAX_URIDA_M3 3
`define AXI_MAX_UWIDA_M3 5
`define AXI_LOG2_MAX_UWIDA_M3 3
`define AXI_RI_LIMIT_M3 0
`define AXI_MAX_RCA_ID_M4 4
`define AXI_LOG2_MAX_RCA_ID_P1_M4 3
`define AXI_MAX_WCA_ID_M4 4
`define AXI_LOG2_MAX_WCA_ID_P1_M4 3
`define AXI_MAX_URIDA_M4 5
`define AXI_LOG2_MAX_URIDA_M4 3
`define AXI_MAX_UWIDA_M4 5
`define AXI_LOG2_MAX_UWIDA_M4 3
`define AXI_RI_LIMIT_M4 0
`define AXI_MAX_RCA_ID_M5 4
`define AXI_LOG2_MAX_RCA_ID_P1_M5 3
`define AXI_MAX_WCA_ID_M5 4
`define AXI_LOG2_MAX_WCA_ID_P1_M5 3
`define AXI_MAX_URIDA_M5 5
`define AXI_LOG2_MAX_URIDA_M5 3
`define AXI_MAX_UWIDA_M5 5
`define AXI_LOG2_MAX_UWIDA_M5 3
`define AXI_RI_LIMIT_M5 0
`define AXI_MAX_RCA_ID_M6 4
`define AXI_LOG2_MAX_RCA_ID_P1_M6 3
`define AXI_MAX_WCA_ID_M6 4
`define AXI_LOG2_MAX_WCA_ID_P1_M6 3
`define AXI_MAX_URIDA_M6 5
`define AXI_LOG2_MAX_URIDA_M6 3
`define AXI_MAX_UWIDA_M6 5
`define AXI_LOG2_MAX_UWIDA_M6 3
`define AXI_RI_LIMIT_M6 0
`define AXI_MAX_RCA_ID_M7 4
`define AXI_LOG2_MAX_RCA_ID_P1_M7 3
`define AXI_MAX_WCA_ID_M7 4
`define AXI_LOG2_MAX_WCA_ID_P1_M7 3
`define AXI_MAX_URIDA_M7 5
`define AXI_LOG2_MAX_URIDA_M7 3
`define AXI_MAX_UWIDA_M7 5
`define AXI_LOG2_MAX_UWIDA_M7 3
`define AXI_RI_LIMIT_M7 0
`define AXI_MAX_RCA_ID_M8 4
`define AXI_LOG2_MAX_RCA_ID_P1_M8 3
`define AXI_MAX_WCA_ID_M8 4
`define AXI_LOG2_MAX_WCA_ID_P1_M8 3
`define AXI_MAX_URIDA_M8 5
`define AXI_LOG2_MAX_URIDA_M8 3
`define AXI_MAX_UWIDA_M8 5
`define AXI_LOG2_MAX_UWIDA_M8 3
`define AXI_RI_LIMIT_M8 0
`define AXI_MAX_RCA_ID_M9 4
`define AXI_LOG2_MAX_RCA_ID_P1_M9 3
`define AXI_MAX_WCA_ID_M9 4
`define AXI_LOG2_MAX_WCA_ID_P1_M9 3
`define AXI_MAX_URIDA_M9 5
`define AXI_LOG2_MAX_URIDA_M9 3
`define AXI_MAX_UWIDA_M9 5
`define AXI_LOG2_MAX_UWIDA_M9 3
`define AXI_RI_LIMIT_M9 0
`define AXI_MAX_RCA_ID_M10 4
`define AXI_LOG2_MAX_RCA_ID_P1_M10 3
`define AXI_MAX_WCA_ID_M10 4
`define AXI_LOG2_MAX_WCA_ID_P1_M10 3
`define AXI_MAX_URIDA_M10 5
`define AXI_LOG2_MAX_URIDA_M10 3
`define AXI_MAX_UWIDA_M10 5
`define AXI_LOG2_MAX_UWIDA_M10 3
`define AXI_RI_LIMIT_M10 0
`define AXI_MAX_RCA_ID_M11 4
`define AXI_LOG2_MAX_RCA_ID_P1_M11 3
`define AXI_MAX_WCA_ID_M11 4
`define AXI_LOG2_MAX_WCA_ID_P1_M11 3
`define AXI_MAX_URIDA_M11 5
`define AXI_LOG2_MAX_URIDA_M11 3
`define AXI_MAX_UWIDA_M11 5
`define AXI_LOG2_MAX_UWIDA_M11 3
`define AXI_RI_LIMIT_M11 0
`define AXI_MAX_RCA_ID_M12 4
`define AXI_LOG2_MAX_RCA_ID_P1_M12 3
`define AXI_MAX_WCA_ID_M12 4
`define AXI_LOG2_MAX_WCA_ID_P1_M12 3
`define AXI_MAX_URIDA_M12 5
`define AXI_LOG2_MAX_URIDA_M12 3
`define AXI_MAX_UWIDA_M12 5
`define AXI_LOG2_MAX_UWIDA_M12 3
`define AXI_RI_LIMIT_M12 0
`define AXI_MAX_RCA_ID_M13 4
`define AXI_LOG2_MAX_RCA_ID_P1_M13 3
`define AXI_MAX_WCA_ID_M13 4
`define AXI_LOG2_MAX_WCA_ID_P1_M13 3
`define AXI_MAX_URIDA_M13 5
`define AXI_LOG2_MAX_URIDA_M13 3
`define AXI_MAX_UWIDA_M13 5
`define AXI_LOG2_MAX_UWIDA_M13 3
`define AXI_RI_LIMIT_M13 0
`define AXI_MAX_RCA_ID_M14 4
`define AXI_LOG2_MAX_RCA_ID_P1_M14 3
`define AXI_MAX_WCA_ID_M14 4
`define AXI_LOG2_MAX_WCA_ID_P1_M14 3
`define AXI_MAX_URIDA_M14 5
`define AXI_LOG2_MAX_URIDA_M14 3
`define AXI_MAX_UWIDA_M14 5
`define AXI_LOG2_MAX_UWIDA_M14 3
`define AXI_RI_LIMIT_M14 0
`define AXI_MAX_RCA_ID_M15 4
`define AXI_LOG2_MAX_RCA_ID_P1_M15 3
`define AXI_MAX_WCA_ID_M15 4
`define AXI_LOG2_MAX_WCA_ID_P1_M15 3
`define AXI_MAX_URIDA_M15 5
`define AXI_LOG2_MAX_URIDA_M15 3
`define AXI_MAX_UWIDA_M15 5
`define AXI_LOG2_MAX_UWIDA_M15 3
`define AXI_RI_LIMIT_M15 0
`define AXI_MAX_RCA_ID_M16 4
`define AXI_LOG2_MAX_RCA_ID_P1_M16 3
`define AXI_MAX_WCA_ID_M16 4
`define AXI_LOG2_MAX_WCA_ID_P1_M16 3
`define AXI_MAX_URIDA_M16 5
`define AXI_LOG2_MAX_URIDA_M16 3
`define AXI_MAX_UWIDA_M16 5
`define AXI_LOG2_MAX_UWIDA_M16 3
`define AXI_RI_LIMIT_M16 0
`define AXI_MAX_FAWC_S0 1
`define AXI_LOG2_MAX_FAWC_S0 1
`define AXI_LOG2_MAX_FAWC_P1_S0 1
`define AXI_MAX_FARC_S0 1
`define AXI_LOG2_MAX_FARC_P1_S0 1
`define AXI_WID_S0 1
`define AXI_MAX_FAC_EN 0
`define AXI_WID_S1 1
`define AXI_LOG2_WID_S1 1
`define AXI_LOG2_WID_P1_S1 1
`define AXI_MAX_FAWC_S1 4
`define AXI_LOG2_MAX_FAWC_S1 2
`define AXI_LOG2_MAX_FAWC_P1_S1 3
`define AXI_MAX_FARC_S1 4
`define AXI_LOG2_MAX_FARC_P1_S1 3
`define AXI_WID_S2 1
`define AXI_LOG2_WID_S2 1
`define AXI_LOG2_WID_P1_S2 1
`define AXI_MAX_FAWC_S2 4
`define AXI_LOG2_MAX_FAWC_S2 2
`define AXI_LOG2_MAX_FAWC_P1_S2 3
`define AXI_MAX_FARC_S2 4
`define AXI_LOG2_MAX_FARC_P1_S2 3
`define AXI_WID_S3 1
`define AXI_LOG2_WID_S3 1
`define AXI_LOG2_WID_P1_S3 1
`define AXI_MAX_FAWC_S3 4
`define AXI_LOG2_MAX_FAWC_S3 2
`define AXI_LOG2_MAX_FAWC_P1_S3 3
`define AXI_MAX_FARC_S3 4
`define AXI_LOG2_MAX_FARC_P1_S3 3
`define AXI_WID_S4 1
`define AXI_LOG2_WID_S4 1
`define AXI_LOG2_WID_P1_S4 1
`define AXI_MAX_FAWC_S4 4
`define AXI_LOG2_MAX_FAWC_S4 2
`define AXI_LOG2_MAX_FAWC_P1_S4 3
`define AXI_MAX_FARC_S4 4
`define AXI_LOG2_MAX_FARC_P1_S4 3
`define AXI_WID_S5 1
`define AXI_LOG2_WID_S5 1
`define AXI_LOG2_WID_P1_S5 1
`define AXI_MAX_FAWC_S5 4
`define AXI_LOG2_MAX_FAWC_S5 2
`define AXI_LOG2_MAX_FAWC_P1_S5 3
`define AXI_MAX_FARC_S5 4
`define AXI_LOG2_MAX_FARC_P1_S5 3
`define AXI_WID_S6 1
`define AXI_LOG2_WID_S6 1
`define AXI_LOG2_WID_P1_S6 1
`define AXI_MAX_FAWC_S6 4
`define AXI_LOG2_MAX_FAWC_S6 2
`define AXI_LOG2_MAX_FAWC_P1_S6 3
`define AXI_MAX_FARC_S6 4
`define AXI_LOG2_MAX_FARC_P1_S6 3
`define AXI_WID_S7 1
`define AXI_LOG2_WID_S7 1
`define AXI_LOG2_WID_P1_S7 1
`define AXI_MAX_FAWC_S7 4
`define AXI_LOG2_MAX_FAWC_S7 2
`define AXI_LOG2_MAX_FAWC_P1_S7 3
`define AXI_MAX_FARC_S7 4
`define AXI_LOG2_MAX_FARC_P1_S7 3
`define AXI_WID_S8 1
`define AXI_LOG2_WID_S8 1
`define AXI_LOG2_WID_P1_S8 1
`define AXI_MAX_FAWC_S8 4
`define AXI_LOG2_MAX_FAWC_S8 2
`define AXI_LOG2_MAX_FAWC_P1_S8 3
`define AXI_MAX_FARC_S8 4
`define AXI_LOG2_MAX_FARC_P1_S8 3
`define AXI_WID_S9 1
`define AXI_LOG2_WID_S9 1
`define AXI_LOG2_WID_P1_S9 1
`define AXI_MAX_FAWC_S9 4
`define AXI_LOG2_MAX_FAWC_S9 2
`define AXI_LOG2_MAX_FAWC_P1_S9 3
`define AXI_MAX_FARC_S9 4
`define AXI_LOG2_MAX_FARC_P1_S9 3
`define AXI_WID_S10 1
`define AXI_LOG2_WID_S10 1
`define AXI_LOG2_WID_P1_S10 1
`define AXI_MAX_FAWC_S10 4
`define AXI_LOG2_MAX_FAWC_S10 2
`define AXI_LOG2_MAX_FAWC_P1_S10 3
`define AXI_MAX_FARC_S10 4
`define AXI_LOG2_MAX_FARC_P1_S10 3
`define AXI_WID_S11 1
`define AXI_LOG2_WID_S11 1
`define AXI_LOG2_WID_P1_S11 1
`define AXI_MAX_FAWC_S11 4
`define AXI_LOG2_MAX_FAWC_S11 2
`define AXI_LOG2_MAX_FAWC_P1_S11 3
`define AXI_MAX_FARC_S11 4
`define AXI_LOG2_MAX_FARC_P1_S11 3
`define AXI_WID_S12 1
`define AXI_LOG2_WID_S12 1
`define AXI_LOG2_WID_P1_S12 1
`define AXI_MAX_FAWC_S12 4
`define AXI_LOG2_MAX_FAWC_S12 2
`define AXI_LOG2_MAX_FAWC_P1_S12 3
`define AXI_MAX_FARC_S12 4
`define AXI_LOG2_MAX_FARC_P1_S12 3
`define AXI_WID_S13 1
`define AXI_LOG2_WID_S13 1
`define AXI_LOG2_WID_P1_S13 1
`define AXI_MAX_FAWC_S13 4
`define AXI_LOG2_MAX_FAWC_S13 2
`define AXI_LOG2_MAX_FAWC_P1_S13 3
`define AXI_MAX_FARC_S13 4
`define AXI_LOG2_MAX_FARC_P1_S13 3
`define AXI_WID_S14 1
`define AXI_LOG2_WID_S14 1
`define AXI_LOG2_WID_P1_S14 1
`define AXI_MAX_FAWC_S14 4
`define AXI_LOG2_MAX_FAWC_S14 2
`define AXI_LOG2_MAX_FAWC_P1_S14 3
`define AXI_MAX_FARC_S14 4
`define AXI_LOG2_MAX_FARC_P1_S14 3
`define AXI_WID_S15 1
`define AXI_LOG2_WID_S15 1
`define AXI_LOG2_WID_P1_S15 1
`define AXI_MAX_FAWC_S15 4
`define AXI_LOG2_MAX_FAWC_S15 2
`define AXI_LOG2_MAX_FAWC_P1_S15 3
`define AXI_MAX_FARC_S15 4
`define AXI_LOG2_MAX_FARC_P1_S15 3
`define AXI_WID_S16 1
`define AXI_LOG2_WID_S16 1
`define AXI_LOG2_WID_P1_S16 1
`define AXI_MAX_FAWC_S16 4
`define AXI_LOG2_MAX_FAWC_S16 2
`define AXI_LOG2_MAX_FAWC_P1_S16 3
`define AXI_MAX_FARC_S16 4
`define AXI_LOG2_MAX_FARC_P1_S16 3
`define AXI_S0_SHARED_FARC 0
`define AXI_LOG2_S0_SHARED_FARC_P1 1
`define AXI_S0_SHARED_AR_HAS_DDCTD 0
`define AXI_S0_SHARED_FAWC 0
`define AXI_LOG2_S0_SHARED_FAWC_P1 1
`define AXI_S0_SHARED_AW_HAS_DDCTD 0
`define AXI_S0_SHARED_W_HAS_DDCTD 0
`define AXI_S1_SHARED_FARC 0
`define AXI_LOG2_S1_SHARED_FARC_P1 1
`define AXI_S1_SHARED_AR_HAS_DDCTD 0
`define AXI_S1_SHARED_FAWC 0
`define AXI_LOG2_S1_SHARED_FAWC_P1 1
`define AXI_S1_SHARED_AW_HAS_DDCTD 0
`define AXI_S1_SHARED_W_HAS_DDCTD 0
`define AXI_S2_SHARED_FARC 0
`define AXI_LOG2_S2_SHARED_FARC_P1 1
`define AXI_S2_SHARED_AR_HAS_DDCTD 0
`define AXI_S2_SHARED_FAWC 0
`define AXI_LOG2_S2_SHARED_FAWC_P1 1
`define AXI_S2_SHARED_AW_HAS_DDCTD 0
`define AXI_S2_SHARED_W_HAS_DDCTD 0
`define AXI_S3_SHARED_FARC 0
`define AXI_LOG2_S3_SHARED_FARC_P1 1
`define AXI_S3_SHARED_AR_HAS_DDCTD 0
`define AXI_S3_SHARED_FAWC 0
`define AXI_LOG2_S3_SHARED_FAWC_P1 1
`define AXI_S3_SHARED_AW_HAS_DDCTD 0
`define AXI_S3_SHARED_W_HAS_DDCTD 0
`define AXI_S4_SHARED_FARC 0
`define AXI_LOG2_S4_SHARED_FARC_P1 1
`define AXI_S4_SHARED_AR_HAS_DDCTD 0
`define AXI_S4_SHARED_FAWC 0
`define AXI_LOG2_S4_SHARED_FAWC_P1 1
`define AXI_S4_SHARED_AW_HAS_DDCTD 0
`define AXI_S4_SHARED_W_HAS_DDCTD 0
`define AXI_S5_SHARED_FARC 0
`define AXI_LOG2_S5_SHARED_FARC_P1 1
`define AXI_S5_SHARED_AR_HAS_DDCTD 0
`define AXI_S5_SHARED_FAWC 0
`define AXI_LOG2_S5_SHARED_FAWC_P1 1
`define AXI_S5_SHARED_AW_HAS_DDCTD 0
`define AXI_S5_SHARED_W_HAS_DDCTD 0
`define AXI_S6_SHARED_FARC 0
`define AXI_LOG2_S6_SHARED_FARC_P1 1
`define AXI_S6_SHARED_AR_HAS_DDCTD 0
`define AXI_S6_SHARED_FAWC 0
`define AXI_LOG2_S6_SHARED_FAWC_P1 1
`define AXI_S6_SHARED_AW_HAS_DDCTD 0
`define AXI_S6_SHARED_W_HAS_DDCTD 0
`define AXI_S7_SHARED_FARC 0
`define AXI_LOG2_S7_SHARED_FARC_P1 1
`define AXI_S7_SHARED_AR_HAS_DDCTD 0
`define AXI_S7_SHARED_FAWC 0
`define AXI_LOG2_S7_SHARED_FAWC_P1 1
`define AXI_S7_SHARED_AW_HAS_DDCTD 0
`define AXI_S7_SHARED_W_HAS_DDCTD 0
`define AXI_S8_SHARED_FARC 0
`define AXI_LOG2_S8_SHARED_FARC_P1 1
`define AXI_S8_SHARED_AR_HAS_DDCTD 0
`define AXI_S8_SHARED_FAWC 0
`define AXI_LOG2_S8_SHARED_FAWC_P1 1
`define AXI_S8_SHARED_AW_HAS_DDCTD 0
`define AXI_S8_SHARED_W_HAS_DDCTD 0
`define AXI_S9_SHARED_FARC 0
`define AXI_LOG2_S9_SHARED_FARC_P1 1
`define AXI_S9_SHARED_AR_HAS_DDCTD 0
`define AXI_S9_SHARED_FAWC 0
`define AXI_LOG2_S9_SHARED_FAWC_P1 1
`define AXI_S9_SHARED_AW_HAS_DDCTD 0
`define AXI_S9_SHARED_W_HAS_DDCTD 0
`define AXI_S10_SHARED_FARC 0
`define AXI_LOG2_S10_SHARED_FARC_P1 1
`define AXI_S10_SHARED_AR_HAS_DDCTD 0
`define AXI_S10_SHARED_FAWC 0
`define AXI_LOG2_S10_SHARED_FAWC_P1 1
`define AXI_S10_SHARED_AW_HAS_DDCTD 0
`define AXI_S10_SHARED_W_HAS_DDCTD 0
`define AXI_S11_SHARED_FARC 0
`define AXI_LOG2_S11_SHARED_FARC_P1 1
`define AXI_S11_SHARED_AR_HAS_DDCTD 0
`define AXI_S11_SHARED_FAWC 0
`define AXI_LOG2_S11_SHARED_FAWC_P1 1
`define AXI_S11_SHARED_AW_HAS_DDCTD 0
`define AXI_S11_SHARED_W_HAS_DDCTD 0
`define AXI_S12_SHARED_FARC 0
`define AXI_LOG2_S12_SHARED_FARC_P1 1
`define AXI_S12_SHARED_AR_HAS_DDCTD 0
`define AXI_S12_SHARED_FAWC 0
`define AXI_LOG2_S12_SHARED_FAWC_P1 1
`define AXI_S12_SHARED_AW_HAS_DDCTD 0
`define AXI_S12_SHARED_W_HAS_DDCTD 0
`define AXI_S13_SHARED_FARC 0
`define AXI_LOG2_S13_SHARED_FARC_P1 1
`define AXI_S13_SHARED_AR_HAS_DDCTD 0
`define AXI_S13_SHARED_FAWC 0
`define AXI_LOG2_S13_SHARED_FAWC_P1 1
`define AXI_S13_SHARED_AW_HAS_DDCTD 0
`define AXI_S13_SHARED_W_HAS_DDCTD 0
`define AXI_S14_SHARED_FARC 0
`define AXI_LOG2_S14_SHARED_FARC_P1 1
`define AXI_S14_SHARED_AR_HAS_DDCTD 0
`define AXI_S14_SHARED_FAWC 0
`define AXI_LOG2_S14_SHARED_FAWC_P1 1
`define AXI_S14_SHARED_AW_HAS_DDCTD 0
`define AXI_S14_SHARED_W_HAS_DDCTD 0
`define AXI_S15_SHARED_FARC 0
`define AXI_LOG2_S15_SHARED_FARC_P1 1
`define AXI_S15_SHARED_AR_HAS_DDCTD 0
`define AXI_S15_SHARED_FAWC 0
`define AXI_LOG2_S15_SHARED_FAWC_P1 1
`define AXI_S15_SHARED_AW_HAS_DDCTD 0
`define AXI_S15_SHARED_W_HAS_DDCTD 0
`define AXI_S16_SHARED_FARC 0
`define AXI_LOG2_S16_SHARED_FARC_P1 1
`define AXI_S16_SHARED_AR_HAS_DDCTD 0
`define AXI_S16_SHARED_FAWC 0
`define AXI_LOG2_S16_SHARED_FAWC_P1 1
`define AXI_S16_SHARED_AW_HAS_DDCTD 0
`define AXI_S16_SHARED_W_HAS_DDCTD 0
`define AXI_M0_SHARED_R_HAS_DDCTD 0
`define AXI_M0_SHARED_B_HAS_DDCTD 0
`define AXI_M1_SHARED_R_HAS_DDCTD 0
`define AXI_M1_SHARED_B_HAS_DDCTD 0
`define AXI_M2_SHARED_R_HAS_DDCTD 0
`define AXI_M2_SHARED_B_HAS_DDCTD 0
`define AXI_M3_SHARED_R_HAS_DDCTD 0
`define AXI_M3_SHARED_B_HAS_DDCTD 0
`define AXI_M4_SHARED_R_HAS_DDCTD 0
`define AXI_M4_SHARED_B_HAS_DDCTD 0
`define AXI_M5_SHARED_R_HAS_DDCTD 0
`define AXI_M5_SHARED_B_HAS_DDCTD 0
`define AXI_M6_SHARED_R_HAS_DDCTD 0
`define AXI_M6_SHARED_B_HAS_DDCTD 0
`define AXI_M7_SHARED_R_HAS_DDCTD 0
`define AXI_M7_SHARED_B_HAS_DDCTD 0
`define AXI_M8_SHARED_R_HAS_DDCTD 0
`define AXI_M8_SHARED_B_HAS_DDCTD 0
`define AXI_M9_SHARED_R_HAS_DDCTD 0
`define AXI_M9_SHARED_B_HAS_DDCTD 0
`define AXI_M10_SHARED_R_HAS_DDCTD 0
`define AXI_M10_SHARED_B_HAS_DDCTD 0
`define AXI_M11_SHARED_R_HAS_DDCTD 0
`define AXI_M11_SHARED_B_HAS_DDCTD 0
`define AXI_M12_SHARED_R_HAS_DDCTD 0
`define AXI_M12_SHARED_B_HAS_DDCTD 0
`define AXI_M13_SHARED_R_HAS_DDCTD 0
`define AXI_M13_SHARED_B_HAS_DDCTD 0
`define AXI_M14_SHARED_R_HAS_DDCTD 0
`define AXI_M14_SHARED_B_HAS_DDCTD 0
`define AXI_M15_SHARED_R_HAS_DDCTD 0
`define AXI_M15_SHARED_B_HAS_DDCTD 0
`define AXI_PRIORITY_M1 0
`define AXI_PRIORITY_M2 0
`define AXI_PRIORITY_M3 0
`define AXI_PRIORITY_M4 0
`define AXI_PRIORITY_M5 0
`define AXI_PRIORITY_M6 0
`define AXI_PRIORITY_M7 0
`define AXI_PRIORITY_M8 0
`define AXI_PRIORITY_M9 0
`define AXI_PRIORITY_M10 0
`define AXI_PRIORITY_M11 0
`define AXI_PRIORITY_M12 0
`define AXI_PRIORITY_M13 0
`define AXI_PRIORITY_M14 0
`define AXI_PRIORITY_M15 0
`define AXI_PRIORITY_M16 0
`define AXI_PRIORITY_S1 1
`define AXI_PRIORITY_S2 1
`define AXI_PRIORITY_S3 1
`define AXI_PRIORITY_S4 1
`define AXI_PRIORITY_S5 1
`define AXI_PRIORITY_S6 1
`define AXI_PRIORITY_S7 1
`define AXI_PRIORITY_S8 1
`define AXI_PRIORITY_S9 1
`define AXI_PRIORITY_S10 1
`define AXI_PRIORITY_S11 1
`define AXI_PRIORITY_S12 1
`define AXI_PRIORITY_S13 1
`define AXI_PRIORITY_S14 1
`define AXI_PRIORITY_S15 1
`define AXI_PRIORITY_S16 1
`define AXI_PRIORITY_S0 0
`define AXI_HAS_EXT_PRIORITY 0
`define AXI_SHARED_LAYER_MASTER_PRIORITY_EN_VAL 0
`define AXI_SHARED_LAYER_MASTER_PRIORITY 1
`define AXI_SHARED_LAYER_SLAVE_PRIORITY_EN_VAL 0
`define AXI_SHARED_LAYER_SLAVE_PRIORITY 1
`define AXI_AR_ARB_TYPE_S0 0
`define AXI_AW_ARB_TYPE_S0 0
`define AXI_AR_ARB_TYPE_S1 0
`define AXI_AW_ARB_TYPE_S1 0
`define AXI_AR_ARB_TYPE_S2 0
`define AXI_AW_ARB_TYPE_S2 0
`define AXI_AR_ARB_TYPE_S3 0
`define AXI_AW_ARB_TYPE_S3 0
`define AXI_AR_ARB_TYPE_S4 0
`define AXI_AW_ARB_TYPE_S4 0
`define AXI_AR_ARB_TYPE_S5 0
`define AXI_AW_ARB_TYPE_S5 0
`define AXI_AR_ARB_TYPE_S6 0
`define AXI_AW_ARB_TYPE_S6 0
`define AXI_AR_ARB_TYPE_S7 0
`define AXI_AW_ARB_TYPE_S7 0
`define AXI_AR_ARB_TYPE_S8 0
`define AXI_AW_ARB_TYPE_S8 0
`define AXI_AR_ARB_TYPE_S9 0
`define AXI_AW_ARB_TYPE_S9 0
`define AXI_AR_ARB_TYPE_S10 0
`define AXI_AW_ARB_TYPE_S10 0
`define AXI_AR_ARB_TYPE_S11 0
`define AXI_AW_ARB_TYPE_S11 0
`define AXI_AR_ARB_TYPE_S12 0
`define AXI_AW_ARB_TYPE_S12 0
`define AXI_AR_ARB_TYPE_S13 0
`define AXI_AW_ARB_TYPE_S13 0
`define AXI_AR_ARB_TYPE_S14 0
`define AXI_AW_ARB_TYPE_S14 0
`define AXI_AR_ARB_TYPE_S15 0
`define AXI_AW_ARB_TYPE_S15 0
`define AXI_AR_ARB_TYPE_S16 0
`define AXI_AW_ARB_TYPE_S16 0
`define AXI_W_ARB_TYPE_S0 0
`define AXI_W_ARB_TYPE_S1 0
`define AXI_W_ARB_TYPE_S2 0
`define AXI_W_ARB_TYPE_S3 0
`define AXI_W_ARB_TYPE_S4 0
`define AXI_W_ARB_TYPE_S5 0
`define AXI_W_ARB_TYPE_S6 0
`define AXI_W_ARB_TYPE_S7 0
`define AXI_W_ARB_TYPE_S8 0
`define AXI_W_ARB_TYPE_S9 0
`define AXI_W_ARB_TYPE_S10 0
`define AXI_W_ARB_TYPE_S11 0
`define AXI_W_ARB_TYPE_S12 0
`define AXI_W_ARB_TYPE_S13 0
`define AXI_W_ARB_TYPE_S14 0
`define AXI_W_ARB_TYPE_S15 0
`define AXI_W_ARB_TYPE_S16 0
`define AXI_R_ARB_TYPE_M1 0
`define AXI_B_ARB_TYPE_M1 0
`define AXI_R_ARB_TYPE_M2 0
`define AXI_B_ARB_TYPE_M2 0
`define AXI_R_ARB_TYPE_M3 0
`define AXI_B_ARB_TYPE_M3 0
`define AXI_R_ARB_TYPE_M4 0
`define AXI_B_ARB_TYPE_M4 0
`define AXI_R_ARB_TYPE_M5 0
`define AXI_B_ARB_TYPE_M5 0
`define AXI_R_ARB_TYPE_M6 0
`define AXI_B_ARB_TYPE_M6 0
`define AXI_R_ARB_TYPE_M7 0
`define AXI_B_ARB_TYPE_M7 0
`define AXI_R_ARB_TYPE_M8 0
`define AXI_B_ARB_TYPE_M8 0
`define AXI_R_ARB_TYPE_M9 0
`define AXI_B_ARB_TYPE_M9 0
`define AXI_R_ARB_TYPE_M10 0
`define AXI_B_ARB_TYPE_M10 0
`define AXI_R_ARB_TYPE_M11 0
`define AXI_B_ARB_TYPE_M11 0
`define AXI_R_ARB_TYPE_M12 0
`define AXI_B_ARB_TYPE_M12 0
`define AXI_R_ARB_TYPE_M13 0
`define AXI_B_ARB_TYPE_M13 0
`define AXI_R_ARB_TYPE_M14 0
`define AXI_B_ARB_TYPE_M14 0
`define AXI_R_ARB_TYPE_M15 0
`define AXI_B_ARB_TYPE_M15 0
`define AXI_R_ARB_TYPE_M16 0
`define AXI_B_ARB_TYPE_M16 0
`define AXI_AR_SHARED_ARB_TYPE 0
`define AXI_AW_SHARED_ARB_TYPE 0
`define AXI_W_SHARED_ARB_TYPE 0
`define AXI_R_SHARED_ARB_TYPE 0
`define AXI_B_SHARED_ARB_TYPE 0
`define AXI_USER_ARB_REMOVAL 1
`define AXI_NUM_RN_S1 1
`define AXI_NUM_RN_S2 1
`define AXI_NUM_RN_S3 1
`define AXI_NUM_RN_S4 1
`define AXI_NUM_RN_S5 1
`define AXI_NUM_RN_S6 1
`define AXI_NUM_RN_S7 1
`define AXI_NUM_RN_S8 1
`define AXI_NUM_RN_S9 1
`define AXI_NUM_RN_S10 1
`define AXI_NUM_RN_S11 1
`define AXI_NUM_RN_S12 1
`define AXI_NUM_RN_S13 1
`define AXI_NUM_RN_S14 1
`define AXI_NUM_RN_S15 1
`define AXI_NUM_RN_S16 1
`define AXI_R1_NSA_S1 32'h60000000
`define AXI_R1_NEA_S1 32'h60000fff
`define AXI_R1_NSA_S2 32'h60001000
`define AXI_R1_NEA_S2 32'h60001fff
`define AXI_R1_NSA_S3 32'h61000000
`define AXI_R1_NEA_S3 32'h61ffffff
`define AXI_R1_NSA_S4 32'he000000
`define AXI_R1_NEA_S4 32'he00ffff
`define AXI_R1_NSA_S5 32'h10000000
`define AXI_R1_NEA_S5 32'h1000ffff
`define AXI_R1_NSA_S6 32'h12000000
`define AXI_R1_NEA_S6 32'h1200ffff
`define AXI_R1_NSA_S7 32'h14000000
`define AXI_R1_NEA_S7 32'h1400ffff
`define AXI_R1_NSA_S8 32'h16000000
`define AXI_R1_NEA_S8 32'h1600ffff
`define AXI_R1_NSA_S9 32'h18000000
`define AXI_R1_NEA_S9 32'h1800ffff
`define AXI_R1_NSA_S10 32'h1a000000
`define AXI_R1_NEA_S10 32'h1a00ffff
`define AXI_R1_NSA_S11 32'h1c000000
`define AXI_R1_NEA_S11 32'h1c00ffff
`define AXI_R1_NSA_S12 32'h1e000000
`define AXI_R1_NEA_S12 32'h1e00ffff
`define AXI_R1_NSA_S13 32'h20000000
`define AXI_R1_NEA_S13 32'h2000ffff
`define AXI_R1_NSA_S14 32'h22000000
`define AXI_R1_NEA_S14 32'h2200ffff
`define AXI_R1_NSA_S15 32'h24000000
`define AXI_R1_NEA_S15 32'h2400ffff
`define AXI_R1_NSA_S16 32'h26000000
`define AXI_R1_NEA_S16 32'h2600ffff
`define AXI_R2_NSA_S1 32'h3000000
`define AXI_R2_NEA_S1 32'h300ffff
`define AXI_R2_NSA_S2 32'hb000000
`define AXI_R2_NEA_S2 32'hb00ffff
`define AXI_R2_NSA_S3 32'hd000000
`define AXI_R2_NEA_S3 32'hd00ffff
`define AXI_R2_NSA_S4 32'hf000000
`define AXI_R2_NEA_S4 32'hf00ffff
`define AXI_R2_NSA_S5 32'h11000000
`define AXI_R2_NEA_S5 32'h1100ffff
`define AXI_R2_NSA_S6 32'h13000000
`define AXI_R2_NEA_S6 32'h1300ffff
`define AXI_R2_NSA_S7 32'h15000000
`define AXI_R2_NEA_S7 32'h1500ffff
`define AXI_R2_NSA_S8 32'h17000000
`define AXI_R2_NEA_S8 32'h1700ffff
`define AXI_R2_NSA_S9 32'h19000000
`define AXI_R2_NEA_S9 32'h1900ffff
`define AXI_R2_NSA_S10 32'h1b000000
`define AXI_R2_NEA_S10 32'h1b00ffff
`define AXI_R2_NSA_S11 32'h1d000000
`define AXI_R2_NEA_S11 32'h1d00ffff
`define AXI_R2_NSA_S12 32'h1f000000
`define AXI_R2_NEA_S12 32'h1f00ffff
`define AXI_R2_NSA_S13 32'h21000000
`define AXI_R2_NEA_S13 32'h2100ffff
`define AXI_R2_NSA_S14 32'h23000000
`define AXI_R2_NEA_S14 32'h2300ffff
`define AXI_R2_NSA_S15 32'h25000000
`define AXI_R2_NEA_S15 32'h2500ffff
`define AXI_R2_NSA_S16 32'h27000000
`define AXI_R2_NEA_S16 32'h2700ffff
`define AXI_R3_NSA_S1 32'h4010000
`define AXI_R3_NEA_S1 32'h401ffff
`define AXI_R3_NSA_S2 32'h4020000
`define AXI_R3_NEA_S2 32'h402ffff
`define AXI_R3_NSA_S3 32'h4030000
`define AXI_R3_NEA_S3 32'h403ffff
`define AXI_R3_NSA_S4 32'h4040000
`define AXI_R3_NEA_S4 32'h404ffff
`define AXI_R3_NSA_S5 32'h4050000
`define AXI_R3_NEA_S5 32'h405ffff
`define AXI_R3_NSA_S6 32'h4060000
`define AXI_R3_NEA_S6 32'h406ffff
`define AXI_R3_NSA_S7 32'h4070000
`define AXI_R3_NEA_S7 32'h407ffff
`define AXI_R3_NSA_S8 32'h4080000
`define AXI_R3_NEA_S8 32'h408ffff
`define AXI_R3_NSA_S9 32'h4090000
`define AXI_R3_NEA_S9 32'h409ffff
`define AXI_R3_NSA_S10 32'h40a0000
`define AXI_R3_NEA_S10 32'h40affff
`define AXI_R3_NSA_S11 32'h40b0000
`define AXI_R3_NEA_S11 32'h40bffff
`define AXI_R3_NSA_S12 32'h40c0000
`define AXI_R3_NEA_S12 32'h40cffff
`define AXI_R3_NSA_S13 32'h40d0000
`define AXI_R3_NEA_S13 32'h40dffff
`define AXI_R3_NSA_S14 32'h40e0000
`define AXI_R3_NEA_S14 32'h40effff
`define AXI_R3_NSA_S15 32'h40f0000
`define AXI_R3_NEA_S15 32'h40fffff
`define AXI_R3_NSA_S16 32'h4000000
`define AXI_R3_NEA_S16 32'h400ffff
`define AXI_R4_NSA_S1 32'h5010000
`define AXI_R4_NEA_S1 32'h501ffff
`define AXI_R4_NSA_S2 32'h5020000
`define AXI_R4_NEA_S2 32'h502ffff
`define AXI_R4_NSA_S3 32'h5030000
`define AXI_R4_NEA_S3 32'h503ffff
`define AXI_R4_NSA_S4 32'h5040000
`define AXI_R4_NEA_S4 32'h504ffff
`define AXI_R4_NSA_S5 32'h5050000
`define AXI_R4_NEA_S5 32'h505ffff
`define AXI_R4_NSA_S6 32'h5060000
`define AXI_R4_NEA_S6 32'h506ffff
`define AXI_R4_NSA_S7 32'h5070000
`define AXI_R4_NEA_S7 32'h507ffff
`define AXI_R4_NSA_S8 32'h5080000
`define AXI_R4_NEA_S8 32'h508ffff
`define AXI_R4_NSA_S9 32'h5090000
`define AXI_R4_NEA_S9 32'h509ffff
`define AXI_R4_NSA_S10 32'h50a0000
`define AXI_R4_NEA_S10 32'h50affff
`define AXI_R4_NSA_S11 32'h50b0000
`define AXI_R4_NEA_S11 32'h50bffff
`define AXI_R4_NSA_S12 32'h50c0000
`define AXI_R4_NEA_S12 32'h50cffff
`define AXI_R4_NSA_S13 32'h50d0000
`define AXI_R4_NEA_S13 32'h50dffff
`define AXI_R4_NSA_S14 32'h50e0000
`define AXI_R4_NEA_S14 32'h50effff
`define AXI_R4_NSA_S15 32'h50f0000
`define AXI_R4_NEA_S15 32'h50fffff
`define AXI_R4_NSA_S16 32'h5000000
`define AXI_R4_NEA_S16 32'h500ffff
`define AXI_R5_NSA_S1 32'h6010000
`define AXI_R5_NEA_S1 32'h601ffff
`define AXI_R5_NSA_S2 32'h6020000
`define AXI_R5_NEA_S2 32'h602ffff
`define AXI_R5_NSA_S3 32'h6030000
`define AXI_R5_NEA_S3 32'h603ffff
`define AXI_R5_NSA_S4 32'h6040000
`define AXI_R5_NEA_S4 32'h604ffff
`define AXI_R5_NSA_S5 32'h6050000
`define AXI_R5_NEA_S5 32'h605ffff
`define AXI_R5_NSA_S6 32'h6060000
`define AXI_R5_NEA_S6 32'h606ffff
`define AXI_R5_NSA_S7 32'h6070000
`define AXI_R5_NEA_S7 32'h607ffff
`define AXI_R5_NSA_S8 32'h6080000
`define AXI_R5_NEA_S8 32'h608ffff
`define AXI_R5_NSA_S9 32'h6090000
`define AXI_R5_NEA_S9 32'h609ffff
`define AXI_R5_NSA_S10 32'h60a0000
`define AXI_R5_NEA_S10 32'h60affff
`define AXI_R5_NSA_S11 32'h60b0000
`define AXI_R5_NEA_S11 32'h60bffff
`define AXI_R5_NSA_S12 32'h60c0000
`define AXI_R5_NEA_S12 32'h60cffff
`define AXI_R5_NSA_S13 32'h60d0000
`define AXI_R5_NEA_S13 32'h60dffff
`define AXI_R5_NSA_S14 32'h60e0000
`define AXI_R5_NEA_S14 32'h60effff
`define AXI_R5_NSA_S15 32'h60f0000
`define AXI_R5_NEA_S15 32'h60fffff
`define AXI_R5_NSA_S16 32'h6000000
`define AXI_R5_NEA_S16 32'h600ffff
`define AXI_R6_NSA_S1 32'h7010000
`define AXI_R6_NEA_S1 32'h701ffff
`define AXI_R6_NSA_S2 32'h7020000
`define AXI_R6_NEA_S2 32'h702ffff
`define AXI_R6_NSA_S3 32'h7030000
`define AXI_R6_NEA_S3 32'h703ffff
`define AXI_R6_NSA_S4 32'h7040000
`define AXI_R6_NEA_S4 32'h704ffff
`define AXI_R6_NSA_S5 32'h7050000
`define AXI_R6_NEA_S5 32'h705ffff
`define AXI_R6_NSA_S6 32'h7060000
`define AXI_R6_NEA_S6 32'h706ffff
`define AXI_R6_NSA_S7 32'h7070000
`define AXI_R6_NEA_S7 32'h707ffff
`define AXI_R6_NSA_S8 32'h7080000
`define AXI_R6_NEA_S8 32'h708ffff
`define AXI_R6_NSA_S9 32'h7090000
`define AXI_R6_NEA_S9 32'h709ffff
`define AXI_R6_NSA_S10 32'h70a0000
`define AXI_R6_NEA_S10 32'h70affff
`define AXI_R6_NSA_S11 32'h70b0000
`define AXI_R6_NEA_S11 32'h70bffff
`define AXI_R6_NSA_S12 32'h70c0000
`define AXI_R6_NEA_S12 32'h70cffff
`define AXI_R6_NSA_S13 32'h70d0000
`define AXI_R6_NEA_S13 32'h70dffff
`define AXI_R6_NSA_S14 32'h70e0000
`define AXI_R6_NEA_S14 32'h70effff
`define AXI_R6_NSA_S15 32'h70f0000
`define AXI_R6_NEA_S15 32'h70fffff
`define AXI_R6_NSA_S16 32'h7000000
`define AXI_R6_NEA_S16 32'h700ffff
`define AXI_R7_NSA_S1 32'h8010000
`define AXI_R7_NEA_S1 32'h801ffff
`define AXI_R7_NSA_S2 32'h8020000
`define AXI_R7_NEA_S2 32'h802ffff
`define AXI_R7_NSA_S3 32'h8030000
`define AXI_R7_NEA_S3 32'h803ffff
`define AXI_R7_NSA_S4 32'h8040000
`define AXI_R7_NEA_S4 32'h804ffff
`define AXI_R7_NSA_S5 32'h8050000
`define AXI_R7_NEA_S5 32'h805ffff
`define AXI_R7_NSA_S6 32'h8060000
`define AXI_R7_NEA_S6 32'h806ffff
`define AXI_R7_NSA_S7 32'h8070000
`define AXI_R7_NEA_S7 32'h807ffff
`define AXI_R7_NSA_S8 32'h8080000
`define AXI_R7_NEA_S8 32'h808ffff
`define AXI_R7_NSA_S9 32'h8090000
`define AXI_R7_NEA_S9 32'h809ffff
`define AXI_R7_NSA_S10 32'h80a0000
`define AXI_R7_NEA_S10 32'h80affff
`define AXI_R7_NSA_S11 32'h80b0000
`define AXI_R7_NEA_S11 32'h80bffff
`define AXI_R7_NSA_S12 32'h80c0000
`define AXI_R7_NEA_S12 32'h80cffff
`define AXI_R7_NSA_S13 32'h80d0000
`define AXI_R7_NEA_S13 32'h80dffff
`define AXI_R7_NSA_S14 32'h80e0000
`define AXI_R7_NEA_S14 32'h80effff
`define AXI_R7_NSA_S15 32'h80f0000
`define AXI_R7_NEA_S15 32'h80fffff
`define AXI_R7_NSA_S16 32'h8000000
`define AXI_R7_NEA_S16 32'h800ffff
`define AXI_R8_NSA_S1 32'h9010000
`define AXI_R8_NEA_S1 32'h901ffff
`define AXI_R8_NSA_S2 32'h9020000
`define AXI_R8_NEA_S2 32'h902ffff
`define AXI_R8_NSA_S3 32'h9030000
`define AXI_R8_NEA_S3 32'h903ffff
`define AXI_R8_NSA_S4 32'h9040000
`define AXI_R8_NEA_S4 32'h904ffff
`define AXI_R8_NSA_S5 32'h9050000
`define AXI_R8_NEA_S5 32'h905ffff
`define AXI_R8_NSA_S6 32'h9060000
`define AXI_R8_NEA_S6 32'h906ffff
`define AXI_R8_NSA_S7 32'h9070000
`define AXI_R8_NEA_S7 32'h907ffff
`define AXI_R8_NSA_S8 32'h9080000
`define AXI_R8_NEA_S8 32'h908ffff
`define AXI_R8_NSA_S9 32'h9090000
`define AXI_R8_NEA_S9 32'h909ffff
`define AXI_R8_NSA_S10 32'h90a0000
`define AXI_R8_NEA_S10 32'h90affff
`define AXI_R8_NSA_S11 32'h90b0000
`define AXI_R8_NEA_S11 32'h90bffff
`define AXI_R8_NSA_S12 32'h90c0000
`define AXI_R8_NEA_S12 32'h90cffff
`define AXI_R8_NSA_S13 32'h90d0000
`define AXI_R8_NEA_S13 32'h90dffff
`define AXI_R8_NSA_S14 32'h90e0000
`define AXI_R8_NEA_S14 32'h90effff
`define AXI_R8_NSA_S15 32'h90f0000
`define AXI_R8_NEA_S15 32'h90fffff
`define AXI_R8_NSA_S16 32'h9000000
`define AXI_R8_NEA_S16 32'h900ffff
`define AXI_NUM_RB_S1 1
`define AXI_NUM_RB_S2 1
`define AXI_NUM_RB_S3 1
`define AXI_NUM_RB_S4 1
`define AXI_NUM_RB_S5 1
`define AXI_NUM_RB_S6 1
`define AXI_NUM_RB_S7 1
`define AXI_NUM_RB_S8 1
`define AXI_NUM_RB_S9 1
`define AXI_NUM_RB_S10 1
`define AXI_NUM_RB_S11 1
`define AXI_NUM_RB_S12 1
`define AXI_NUM_RB_S13 1
`define AXI_NUM_RB_S14 1
`define AXI_NUM_RB_S15 1
`define AXI_NUM_RB_S16 1
`define AXI_R1_BSA_S1 32'h60000000
`define AXI_R1_BEA_S1 32'h60000fff
`define AXI_R1_BSA_S2 32'h60001000
`define AXI_R1_BEA_S2 32'h60001fff
`define AXI_R1_BSA_S3 32'h61000000
`define AXI_R1_BEA_S3 32'h61ffffff
`define AXI_R1_BSA_S4 32'he000000
`define AXI_R1_BEA_S4 32'he00ffff
`define AXI_R1_BSA_S5 32'h10000000
`define AXI_R1_BEA_S5 32'h1000ffff
`define AXI_R1_BSA_S6 32'h12000000
`define AXI_R1_BEA_S6 32'h1200ffff
`define AXI_R1_BSA_S7 32'h14000000
`define AXI_R1_BEA_S7 32'h1400ffff
`define AXI_R1_BSA_S8 32'h16000000
`define AXI_R1_BEA_S8 32'h1600ffff
`define AXI_R1_BSA_S9 32'h18000000
`define AXI_R1_BEA_S9 32'h1800ffff
`define AXI_R1_BSA_S10 32'h1a000000
`define AXI_R1_BEA_S10 32'h1a00ffff
`define AXI_R1_BSA_S11 32'h1c000000
`define AXI_R1_BEA_S11 32'h1c00ffff
`define AXI_R1_BSA_S12 32'h1e000000
`define AXI_R1_BEA_S12 32'h1e00ffff
`define AXI_R1_BSA_S13 32'h20000000
`define AXI_R1_BEA_S13 32'h2000ffff
`define AXI_R1_BSA_S14 32'h22000000
`define AXI_R1_BEA_S14 32'h2200ffff
`define AXI_R1_BSA_S15 32'h24000000
`define AXI_R1_BEA_S15 32'h2400ffff
`define AXI_R1_BSA_S16 32'h26000000
`define AXI_R1_BEA_S16 32'h2600ffff
`define AXI_R2_BSA_S1 32'h3000000
`define AXI_R2_BEA_S1 32'h300ffff
`define AXI_R2_BSA_S2 32'hb000000
`define AXI_R2_BEA_S2 32'hb00ffff
`define AXI_R2_BSA_S3 32'hd000000
`define AXI_R2_BEA_S3 32'hd00ffff
`define AXI_R2_BSA_S4 32'hf000000
`define AXI_R2_BEA_S4 32'hf00ffff
`define AXI_R2_BSA_S5 32'h11000000
`define AXI_R2_BEA_S5 32'h1100ffff
`define AXI_R2_BSA_S6 32'h13000000
`define AXI_R2_BEA_S6 32'h1300ffff
`define AXI_R2_BSA_S7 32'h15000000
`define AXI_R2_BEA_S7 32'h1500ffff
`define AXI_R2_BSA_S8 32'h17000000
`define AXI_R2_BEA_S8 32'h1700ffff
`define AXI_R2_BSA_S9 32'h19000000
`define AXI_R2_BEA_S9 32'h1900ffff
`define AXI_R2_BSA_S10 32'h1b000000
`define AXI_R2_BEA_S10 32'h1b00ffff
`define AXI_R2_BSA_S11 32'h1d000000
`define AXI_R2_BEA_S11 32'h1d00ffff
`define AXI_R2_BSA_S12 32'h1f000000
`define AXI_R2_BEA_S12 32'h1f00ffff
`define AXI_R2_BSA_S13 32'h21000000
`define AXI_R2_BEA_S13 32'h2100ffff
`define AXI_R2_BSA_S14 32'h23000000
`define AXI_R2_BEA_S14 32'h2300ffff
`define AXI_R2_BSA_S15 32'h25000000
`define AXI_R2_BEA_S15 32'h2500ffff
`define AXI_R2_BSA_S16 32'h27000000
`define AXI_R2_BEA_S16 32'h2700ffff
`define AXI_R3_BSA_S1 32'h4010000
`define AXI_R3_BEA_S1 32'h401ffff
`define AXI_R3_BSA_S2 32'h4020000
`define AXI_R3_BEA_S2 32'h402ffff
`define AXI_R3_BSA_S3 32'h4030000
`define AXI_R3_BEA_S3 32'h403ffff
`define AXI_R3_BSA_S4 32'h4040000
`define AXI_R3_BEA_S4 32'h404ffff
`define AXI_R3_BSA_S5 32'h4050000
`define AXI_R3_BEA_S5 32'h405ffff
`define AXI_R3_BSA_S6 32'h4060000
`define AXI_R3_BEA_S6 32'h406ffff
`define AXI_R3_BSA_S7 32'h4070000
`define AXI_R3_BEA_S7 32'h407ffff
`define AXI_R3_BSA_S8 32'h4080000
`define AXI_R3_BEA_S8 32'h408ffff
`define AXI_R3_BSA_S9 32'h4090000
`define AXI_R3_BEA_S9 32'h409ffff
`define AXI_R3_BSA_S10 32'h40a0000
`define AXI_R3_BEA_S10 32'h40affff
`define AXI_R3_BSA_S11 32'h40b0000
`define AXI_R3_BEA_S11 32'h40bffff
`define AXI_R3_BSA_S12 32'h40c0000
`define AXI_R3_BEA_S12 32'h40cffff
`define AXI_R3_BSA_S13 32'h40d0000
`define AXI_R3_BEA_S13 32'h40dffff
`define AXI_R3_BSA_S14 32'h40e0000
`define AXI_R3_BEA_S14 32'h40effff
`define AXI_R3_BSA_S15 32'h40f0000
`define AXI_R3_BEA_S15 32'h40fffff
`define AXI_R3_BSA_S16 32'h4000000
`define AXI_R3_BEA_S16 32'h400ffff
`define AXI_R4_BSA_S1 32'h5010000
`define AXI_R4_BEA_S1 32'h501ffff
`define AXI_R4_BSA_S2 32'h5020000
`define AXI_R4_BEA_S2 32'h502ffff
`define AXI_R4_BSA_S3 32'h5030000
`define AXI_R4_BEA_S3 32'h503ffff
`define AXI_R4_BSA_S4 32'h5040000
`define AXI_R4_BEA_S4 32'h504ffff
`define AXI_R4_BSA_S5 32'h5050000
`define AXI_R4_BEA_S5 32'h505ffff
`define AXI_R4_BSA_S6 32'h5060000
`define AXI_R4_BEA_S6 32'h506ffff
`define AXI_R4_BSA_S7 32'h5070000
`define AXI_R4_BEA_S7 32'h507ffff
`define AXI_R4_BSA_S8 32'h5080000
`define AXI_R4_BEA_S8 32'h508ffff
`define AXI_R4_BSA_S9 32'h5090000
`define AXI_R4_BEA_S9 32'h509ffff
`define AXI_R4_BSA_S10 32'h50a0000
`define AXI_R4_BEA_S10 32'h50affff
`define AXI_R4_BSA_S11 32'h50b0000
`define AXI_R4_BEA_S11 32'h50bffff
`define AXI_R4_BSA_S12 32'h50c0000
`define AXI_R4_BEA_S12 32'h50cffff
`define AXI_R4_BSA_S13 32'h50d0000
`define AXI_R4_BEA_S13 32'h50dffff
`define AXI_R4_BSA_S14 32'h50e0000
`define AXI_R4_BEA_S14 32'h50effff
`define AXI_R4_BSA_S15 32'h50f0000
`define AXI_R4_BEA_S15 32'h50fffff
`define AXI_R4_BSA_S16 32'h5000000
`define AXI_R4_BEA_S16 32'h500ffff
`define AXI_R5_BSA_S1 32'h6010000
`define AXI_R5_BEA_S1 32'h601ffff
`define AXI_R5_BSA_S2 32'h6020000
`define AXI_R5_BEA_S2 32'h602ffff
`define AXI_R5_BSA_S3 32'h6030000
`define AXI_R5_BEA_S3 32'h603ffff
`define AXI_R5_BSA_S4 32'h6040000
`define AXI_R5_BEA_S4 32'h604ffff
`define AXI_R5_BSA_S5 32'h6050000
`define AXI_R5_BEA_S5 32'h605ffff
`define AXI_R5_BSA_S6 32'h6060000
`define AXI_R5_BEA_S6 32'h606ffff
`define AXI_R5_BSA_S7 32'h6070000
`define AXI_R5_BEA_S7 32'h607ffff
`define AXI_R5_BSA_S8 32'h6080000
`define AXI_R5_BEA_S8 32'h608ffff
`define AXI_R5_BSA_S9 32'h6090000
`define AXI_R5_BEA_S9 32'h609ffff
`define AXI_R5_BSA_S10 32'h60a0000
`define AXI_R5_BEA_S10 32'h60affff
`define AXI_R5_BSA_S11 32'h60b0000
`define AXI_R5_BEA_S11 32'h60bffff
`define AXI_R5_BSA_S12 32'h60c0000
`define AXI_R5_BEA_S12 32'h60cffff
`define AXI_R5_BSA_S13 32'h60d0000
`define AXI_R5_BEA_S13 32'h60dffff
`define AXI_R5_BSA_S14 32'h60e0000
`define AXI_R5_BEA_S14 32'h60effff
`define AXI_R5_BSA_S15 32'h60f0000
`define AXI_R5_BEA_S15 32'h60fffff
`define AXI_R5_BSA_S16 32'h6000000
`define AXI_R5_BEA_S16 32'h600ffff
`define AXI_R6_BSA_S1 32'h7010000
`define AXI_R6_BEA_S1 32'h701ffff
`define AXI_R6_BSA_S2 32'h7020000
`define AXI_R6_BEA_S2 32'h702ffff
`define AXI_R6_BSA_S3 32'h7030000
`define AXI_R6_BEA_S3 32'h703ffff
`define AXI_R6_BSA_S4 32'h7040000
`define AXI_R6_BEA_S4 32'h704ffff
`define AXI_R6_BSA_S5 32'h7050000
`define AXI_R6_BEA_S5 32'h705ffff
`define AXI_R6_BSA_S6 32'h7060000
`define AXI_R6_BEA_S6 32'h706ffff
`define AXI_R6_BSA_S7 32'h7070000
`define AXI_R6_BEA_S7 32'h707ffff
`define AXI_R6_BSA_S8 32'h7080000
`define AXI_R6_BEA_S8 32'h708ffff
`define AXI_R6_BSA_S9 32'h7090000
`define AXI_R6_BEA_S9 32'h709ffff
`define AXI_R6_BSA_S10 32'h70a0000
`define AXI_R6_BEA_S10 32'h70affff
`define AXI_R6_BSA_S11 32'h70b0000
`define AXI_R6_BEA_S11 32'h70bffff
`define AXI_R6_BSA_S12 32'h70c0000
`define AXI_R6_BEA_S12 32'h70cffff
`define AXI_R6_BSA_S13 32'h70d0000
`define AXI_R6_BEA_S13 32'h70dffff
`define AXI_R6_BSA_S14 32'h70e0000
`define AXI_R6_BEA_S14 32'h70effff
`define AXI_R6_BSA_S15 32'h70f0000
`define AXI_R6_BEA_S15 32'h70fffff
`define AXI_R6_BSA_S16 32'h7000000
`define AXI_R6_BEA_S16 32'h700ffff
`define AXI_R7_BSA_S1 32'h8010000
`define AXI_R7_BEA_S1 32'h801ffff
`define AXI_R7_BSA_S2 32'h8020000
`define AXI_R7_BEA_S2 32'h802ffff
`define AXI_R7_BSA_S3 32'h8030000
`define AXI_R7_BEA_S3 32'h803ffff
`define AXI_R7_BSA_S4 32'h8040000
`define AXI_R7_BEA_S4 32'h804ffff
`define AXI_R7_BSA_S5 32'h8050000
`define AXI_R7_BEA_S5 32'h805ffff
`define AXI_R7_BSA_S6 32'h8060000
`define AXI_R7_BEA_S6 32'h806ffff
`define AXI_R7_BSA_S7 32'h8070000
`define AXI_R7_BEA_S7 32'h807ffff
`define AXI_R7_BSA_S8 32'h8080000
`define AXI_R7_BEA_S8 32'h808ffff
`define AXI_R7_BSA_S9 32'h8090000
`define AXI_R7_BEA_S9 32'h809ffff
`define AXI_R7_BSA_S10 32'h80a0000
`define AXI_R7_BEA_S10 32'h80affff
`define AXI_R7_BSA_S11 32'h80b0000
`define AXI_R7_BEA_S11 32'h80bffff
`define AXI_R7_BSA_S12 32'h80c0000
`define AXI_R7_BEA_S12 32'h80cffff
`define AXI_R7_BSA_S13 32'h80d0000
`define AXI_R7_BEA_S13 32'h80dffff
`define AXI_R7_BSA_S14 32'h80e0000
`define AXI_R7_BEA_S14 32'h80effff
`define AXI_R7_BSA_S15 32'h80f0000
`define AXI_R7_BEA_S15 32'h80fffff
`define AXI_R7_BSA_S16 32'h8000000
`define AXI_R7_BEA_S16 32'h800ffff
`define AXI_R8_BSA_S1 32'h9010000
`define AXI_R8_BEA_S1 32'h901ffff
`define AXI_R8_BSA_S2 32'h9020000
`define AXI_R8_BEA_S2 32'h902ffff
`define AXI_R8_BSA_S3 32'h9030000
`define AXI_R8_BEA_S3 32'h903ffff
`define AXI_R8_BSA_S4 32'h9040000
`define AXI_R8_BEA_S4 32'h904ffff
`define AXI_R8_BSA_S5 32'h9050000
`define AXI_R8_BEA_S5 32'h905ffff
`define AXI_R8_BSA_S6 32'h9060000
`define AXI_R8_BEA_S6 32'h906ffff
`define AXI_R8_BSA_S7 32'h9070000
`define AXI_R8_BEA_S7 32'h907ffff
`define AXI_R8_BSA_S8 32'h9080000
`define AXI_R8_BEA_S8 32'h908ffff
`define AXI_R8_BSA_S9 32'h9090000
`define AXI_R8_BEA_S9 32'h909ffff
`define AXI_R8_BSA_S10 32'h90a0000
`define AXI_R8_BEA_S10 32'h90affff
`define AXI_R8_BSA_S11 32'h90b0000
`define AXI_R8_BEA_S11 32'h90bffff
`define AXI_R8_BSA_S12 32'h90c0000
`define AXI_R8_BEA_S12 32'h90cffff
`define AXI_R8_BSA_S13 32'h90d0000
`define AXI_R8_BEA_S13 32'h90dffff
`define AXI_R8_BSA_S14 32'h90e0000
`define AXI_R8_BEA_S14 32'h90effff
`define AXI_R8_BSA_S15 32'h90f0000
`define AXI_R8_BEA_S15 32'h90fffff
`define AXI_R8_BSA_S16 32'h9000000
`define AXI_R8_BEA_S16 32'h900ffff
`define AXI_AR_PYLD_M_W 58
`define AXI_AW_PYLD_M_W 58
`define AXI_W_PYLD_M_W 78
`define AXI_R_PYLD_M_W 72
`define AXI_B_PYLD_M_W 7
`define AXI_AR_PYLD_S_W 59
`define AXI_AW_PYLD_S_W 59
`define AXI_W_PYLD_S_W 79
`define AXI_R_PYLD_S_W 73
`define AXI_B_PYLD_S_W 8
`define AXI_HAS_S0
`define AXI_HAS_S1
`define AXI_HAS_S2
`define AXI_HAS_S3
`define AXI_HAS_M1
`define AXI_HAS_M2
`define AXI_NMV_S0 `AXI_NUM_MASTERS
`define AXI_SYS_NUM_FOR_M1 1
`define AXI_SYS_NUM_FOR_M2 2
`define AXI_SYS_NUM_FOR_M3 3
`define AXI_SYS_NUM_FOR_M4 4
`define AXI_SYS_NUM_FOR_M5 5
`define AXI_SYS_NUM_FOR_M6 6
`define AXI_SYS_NUM_FOR_M7 7
`define AXI_SYS_NUM_FOR_M8 8
`define AXI_SYS_NUM_FOR_M9 9
`define AXI_SYS_NUM_FOR_M10 10
`define AXI_SYS_NUM_FOR_M11 11
`define AXI_SYS_NUM_FOR_M12 12
`define AXI_SYS_NUM_FOR_M13 13
`define AXI_SYS_NUM_FOR_M14 14
`define AXI_SYS_NUM_FOR_M15 15
`define AXI_SYS_NUM_FOR_M16 16
`define AXI_NUM_ICM 0
`define AXI_ACC_NON_LCL_SLV_S1 0
`define AXI_ACC_NON_LCL_SLV_S2 0
`define AXI_ACC_NON_LCL_SLV_S3 0
`define AXI_ACC_NON_LCL_SLV_S4 0
`define AXI_ACC_NON_LCL_SLV_S5 0
`define AXI_ACC_NON_LCL_SLV_S6 0
`define AXI_ACC_NON_LCL_SLV_S7 0
`define AXI_ACC_NON_LCL_SLV_S8 0
`define AXI_ACC_NON_LCL_SLV_S9 0
`define AXI_ACC_NON_LCL_SLV_S10 0
`define AXI_ACC_NON_LCL_SLV_S11 0
`define AXI_ACC_NON_LCL_SLV_S12 0
`define AXI_ACC_NON_LCL_SLV_S13 0
`define AXI_ACC_NON_LCL_SLV_S14 0
`define AXI_ACC_NON_LCL_SLV_S15 0
`define AXI_ACC_NON_LCL_SLV_S16 0
`define AXI_IS_ICM_M1 0
`define AXI_IS_ICM_M2 0
`define AXI_IS_ICM_M3 0
`define AXI_IS_ICM_M4 0
`define AXI_IS_ICM_M5 0
`define AXI_IS_ICM_M6 0
`define AXI_IS_ICM_M7 0
`define AXI_IS_ICM_M8 0
`define AXI_IS_ICM_M9 0
`define AXI_IS_ICM_M10 0
`define AXI_IS_ICM_M11 0
`define AXI_IS_ICM_M12 0
`define AXI_IS_ICM_M13 0
`define AXI_IS_ICM_M14 0
`define AXI_IS_ICM_M15 0
`define AXI_IS_ICM_M16 0
`define AXI_IDW_M1 5
`define AXI_IDW_M2 5
`define AXI_IDW_M3 5
`define AXI_IDW_M4 5
`define AXI_NUM_MST_THRU_ICM1 1
`define AXI_NUM_MST_THRU_ICM2 1
`define AXI_NUM_MST_THRU_ICM3 1
`define AXI_NUM_MST_THRU_ICM4 1
`define AXI_ALLOW_MST1_ICM1 1
`define AXI_ALLOW_MST2_ICM1 1
`define AXI_ALLOW_MST3_ICM1 1
`define AXI_ALLOW_MST4_ICM1 1
`define AXI_ALLOW_MST5_ICM1 1
`define AXI_ALLOW_MST6_ICM1 1
`define AXI_ALLOW_MST7_ICM1 1
`define AXI_ALLOW_MST8_ICM1 1
`define AXI_ALLOW_MST1_ICM2 1
`define AXI_ALLOW_MST2_ICM2 1
`define AXI_ALLOW_MST3_ICM2 1
`define AXI_ALLOW_MST4_ICM2 1
`define AXI_ALLOW_MST5_ICM2 1
`define AXI_ALLOW_MST6_ICM2 1
`define AXI_ALLOW_MST7_ICM2 1
`define AXI_ALLOW_MST8_ICM2 1
`define AXI_ALLOW_MST1_ICM3 1
`define AXI_ALLOW_MST2_ICM3 1
`define AXI_ALLOW_MST3_ICM3 1
`define AXI_ALLOW_MST4_ICM3 1
`define AXI_ALLOW_MST5_ICM3 1
`define AXI_ALLOW_MST6_ICM3 1
`define AXI_ALLOW_MST7_ICM3 1
`define AXI_ALLOW_MST8_ICM3 1
`define AXI_ALLOW_MST1_ICM4 1
`define AXI_ALLOW_MST2_ICM4 1
`define AXI_ALLOW_MST3_ICM4 1
`define AXI_ALLOW_MST4_ICM4 1
`define AXI_ALLOW_MST5_ICM4 1
`define AXI_ALLOW_MST6_ICM4 1
`define AXI_ALLOW_MST7_ICM4 1
`define AXI_ALLOW_MST8_ICM4 1
`define AXI_PNUM_FOR_SYS_NUM_M1 1
`define AXI_PNUM_FOR_SYS_NUM_M2 2
`define AXI_PNUM_FOR_SYS_NUM_M3 0
`define AXI_PNUM_FOR_SYS_NUM_M4 0
`define AXI_PNUM_FOR_SYS_NUM_M5 0
`define AXI_PNUM_FOR_SYS_NUM_M6 0
`define AXI_PNUM_FOR_SYS_NUM_M7 0
`define AXI_PNUM_FOR_SYS_NUM_M8 0
`define AXI_PNUM_FOR_SYS_NUM_M9 0
`define AXI_PNUM_FOR_SYS_NUM_M10 0
`define AXI_PNUM_FOR_SYS_NUM_M11 0
`define AXI_PNUM_FOR_SYS_NUM_M12 0
`define AXI_PNUM_FOR_SYS_NUM_M13 0
`define AXI_PNUM_FOR_SYS_NUM_M14 0
`define AXI_PNUM_FOR_SYS_NUM_M15 0
`define AXI_PNUM_FOR_SYS_NUM_M16 0
`define AXI_PNUM_FOR_SYS_NUM_M17 0
`define AXI_PNUM_FOR_SYS_NUM_M18 0
`define AXI_PNUM_FOR_SYS_NUM_M19 0
`define AXI_PNUM_FOR_SYS_NUM_M20 0
`define AXI_PNUM_FOR_SYS_NUM_M21 0
`define AXI_PNUM_FOR_SYS_NUM_M22 0
`define AXI_PNUM_FOR_SYS_NUM_M23 0
`define AXI_PNUM_FOR_SYS_NUM_M24 0
`define AXI_PNUM_FOR_SYS_NUM_M25 0
`define AXI_PNUM_FOR_SYS_NUM_M26 0
`define AXI_PNUM_FOR_SYS_NUM_M27 0
`define AXI_PNUM_FOR_SYS_NUM_M28 0
`define AXI_PNUM_FOR_SYS_NUM_M29 0
`define AXI_PNUM_FOR_SYS_NUM_M30 0
`define AXI_PNUM_FOR_SYS_NUM_M31 0
`define AXI_PNUM_FOR_SYS_NUM_M32 0
`define AXI_PNUM_FOR_SYS_NUM_M33 0
`define AXI_PNUM_FOR_SYS_NUM_M34 0
`define AXI_PNUM_FOR_SYS_NUM_M35 0
`define AXI_PNUM_FOR_SYS_NUM_M36 0
`define AXI_PNUM_FOR_SYS_NUM_M37 0
`define AXI_PNUM_FOR_SYS_NUM_M38 0
`define AXI_PNUM_FOR_SYS_NUM_M39 0
`define AXI_PNUM_FOR_SYS_NUM_M40 0
`define AXI_PNUM_FOR_SYS_NUM_M41 0
`define AXI_PNUM_FOR_SYS_NUM_M42 0
`define AXI_PNUM_FOR_SYS_NUM_M43 0
`define AXI_PNUM_FOR_SYS_NUM_M44 0
`define AXI_PNUM_FOR_SYS_NUM_M45 0
`define AXI_PNUM_FOR_SYS_NUM_M46 0
`define AXI_PNUM_FOR_SYS_NUM_M47 0
`define AXI_PNUM_FOR_SYS_NUM_M48 0
`define AXI_PNUM_FOR_SYS_NUM_M49 0
`define AXI_PNUM_FOR_SYS_NUM_M50 0
`define AXI_PNUM_FOR_SYS_NUM_M51 0
`define AXI_PNUM_FOR_SYS_NUM_M52 0
`define AXI_PNUM_FOR_SYS_NUM_M53 0
`define AXI_PNUM_FOR_SYS_NUM_M54 0
`define AXI_PNUM_FOR_SYS_NUM_M55 0
`define AXI_PNUM_FOR_SYS_NUM_M56 0
`define AXI_PNUM_FOR_SYS_NUM_M57 0
`define AXI_PNUM_FOR_SYS_NUM_M58 0
`define AXI_PNUM_FOR_SYS_NUM_M59 0
`define AXI_PNUM_FOR_SYS_NUM_M60 0
`define AXI_PNUM_FOR_SYS_NUM_M61 0
`define AXI_PNUM_FOR_SYS_NUM_M62 0
`define AXI_PNUM_FOR_SYS_NUM_M63 0
`define AXI_PNUM_FOR_SYS_NUM_M64 0
`define AXI_SRC_LICENSE_CHK 1
`define AXI_NSPV_M1_AR_QOSARB 0
`define AXI_NSPV_M2_AR_QOSARB 0
`define AXI_NSPV_M3_AR_QOSARB 1
`define AXI_NSPV_M4_AR_QOSARB 1
`define AXI_NSPV_M5_AR_QOSARB 1
`define AXI_NSPV_M6_AR_QOSARB 1
`define AXI_NSPV_M7_AR_QOSARB 1
`define AXI_NSPV_M8_AR_QOSARB 1
`define AXI_NSPV_M9_AR_QOSARB 1
`define AXI_NSPV_M10_AR_QOSARB 1
`define AXI_NSPV_M11_AR_QOSARB 1
`define AXI_NSPV_M12_AR_QOSARB 1
`define AXI_NSPV_M13_AR_QOSARB 1
`define AXI_NSPV_M14_AR_QOSARB 1
`define AXI_NSPV_M15_AR_QOSARB 1
`define AXI_NSPV_M16_AR_QOSARB 1
`define AXI_NSPV_M1_AW_QOSARB 0
`define AXI_NSPV_M2_AW_QOSARB 0
`define AXI_NSPV_M3_AW_QOSARB 1
`define AXI_NSPV_M4_AW_QOSARB 1
`define AXI_NSPV_M5_AW_QOSARB 1
`define AXI_NSPV_M6_AW_QOSARB 1
`define AXI_NSPV_M7_AW_QOSARB 1
`define AXI_NSPV_M8_AW_QOSARB 1
`define AXI_NSPV_M9_AW_QOSARB 1
`define AXI_NSPV_M10_AW_QOSARB 1
`define AXI_NSPV_M11_AW_QOSARB 1
`define AXI_NSPV_M12_AW_QOSARB 1
`define AXI_NSPV_M13_AW_QOSARB 1
`define AXI_NSPV_M14_AW_QOSARB 1
`define AXI_NSPV_M15_AW_QOSARB 1
`define AXI_NSPV_M16_AW_QOSARB 1
`define AXI_AR_HAS_QOS_REGULATOR_M1 0
`define AXI_AR_HAS_QOS_REGULATOR_M2 0
`define AXI_AR_HAS_QOS_REGULATOR_M3 0
`define AXI_AR_HAS_QOS_REGULATOR_M4 0
`define AXI_AR_HAS_QOS_REGULATOR_M5 0
`define AXI_AR_HAS_QOS_REGULATOR_M6 0
`define AXI_AR_HAS_QOS_REGULATOR_M7 0
`define AXI_AR_HAS_QOS_REGULATOR_M8 0
`define AXI_AR_HAS_QOS_REGULATOR_M9 0
`define AXI_AR_HAS_QOS_REGULATOR_M10 0
`define AXI_AR_HAS_QOS_REGULATOR_M11 0
`define AXI_AR_HAS_QOS_REGULATOR_M12 0
`define AXI_AR_HAS_QOS_REGULATOR_M13 0
`define AXI_AR_HAS_QOS_REGULATOR_M14 0
`define AXI_AR_HAS_QOS_REGULATOR_M15 0
`define AXI_AR_HAS_QOS_REGULATOR_M16 0
`define AXI_AW_HAS_QOS_REGULATOR_M1 0
`define AXI_AW_HAS_QOS_REGULATOR_M2 0
`define AXI_AW_HAS_QOS_REGULATOR_M3 0
`define AXI_AW_HAS_QOS_REGULATOR_M4 0
`define AXI_AW_HAS_QOS_REGULATOR_M5 0
`define AXI_AW_HAS_QOS_REGULATOR_M6 0
`define AXI_AW_HAS_QOS_REGULATOR_M7 0
`define AXI_AW_HAS_QOS_REGULATOR_M8 0
`define AXI_AW_HAS_QOS_REGULATOR_M9 0
`define AXI_AW_HAS_QOS_REGULATOR_M10 0
`define AXI_AW_HAS_QOS_REGULATOR_M11 0
`define AXI_AW_HAS_QOS_REGULATOR_M12 0
`define AXI_AW_HAS_QOS_REGULATOR_M13 0
`define AXI_AW_HAS_QOS_REGULATOR_M14 0
`define AXI_AW_HAS_QOS_REGULATOR_M15 0
`define AXI_AW_HAS_QOS_REGULATOR_M16 0
`define AXI_HAS_ARQOS_EXT_M1 0
`define AXI_ARQOS_INT_M1
`define AXI_HAS_ARQOS_EXT_M2 0
`define AXI_ARQOS_INT_M2
`define AXI_HAS_ARQOS_EXT_M3 0
`define AXI_HAS_ARQOS_EXT_M4 0
`define AXI_HAS_ARQOS_EXT_M5 0
`define AXI_HAS_ARQOS_EXT_M6 0
`define AXI_HAS_ARQOS_EXT_M7 0
`define AXI_HAS_ARQOS_EXT_M8 0
`define AXI_HAS_ARQOS_EXT_M9 0
`define AXI_HAS_ARQOS_EXT_M10 0
`define AXI_HAS_ARQOS_EXT_M11 0
`define AXI_HAS_ARQOS_EXT_M12 0
`define AXI_HAS_ARQOS_EXT_M13 0
`define AXI_HAS_ARQOS_EXT_M14 0
`define AXI_HAS_ARQOS_EXT_M15 0
`define AXI_HAS_ARQOS_EXT_M16 0
`define AXI_HAS_AWQOS_EXT_M1 0
`define AXI_AWQOS_INT_M1
`define AXI_HAS_AWQOS_EXT_M2 0
`define AXI_AWQOS_INT_M2
`define AXI_HAS_AWQOS_EXT_M3 0
`define AXI_HAS_AWQOS_EXT_M4 0
`define AXI_HAS_AWQOS_EXT_M5 0
`define AXI_HAS_AWQOS_EXT_M6 0
`define AXI_HAS_AWQOS_EXT_M7 0
`define AXI_HAS_AWQOS_EXT_M8 0
`define AXI_HAS_AWQOS_EXT_M9 0
`define AXI_HAS_AWQOS_EXT_M10 0
`define AXI_HAS_AWQOS_EXT_M11 0
`define AXI_HAS_AWQOS_EXT_M12 0
`define AXI_HAS_AWQOS_EXT_M13 0
`define AXI_HAS_AWQOS_EXT_M14 0
`define AXI_HAS_AWQOS_EXT_M15 0
`define AXI_HAS_AWQOS_EXT_M16 0
`define SNPS_RCE_INTERNAL_ON 
`define AXI_HAS_APB 0
`define AXI_HAS_APB3 0
`define APB_DATA_WIDTH 32
`define AXI_IC_REG_BASE_ADDR 32'h00400
`define AXI_NUM_SYNC_FF 2
`define DW_AXI_VERSION_ID 32'h3430362a
`define AXI_VERIF_EN 1
`define AXI_4 1
`define AXI_ACELITE 0
`define AXI_HAS_REGIONS_S1 0
`define AXI_HAS_REGIONS_S2 0
`define AXI_HAS_REGIONS_S3 0
`define AXI_HAS_REGIONS_S4 0
`define AXI_HAS_REGIONS_S5 0
`define AXI_HAS_REGIONS_S6 0
`define AXI_HAS_REGIONS_S7 0
`define AXI_HAS_REGIONS_S8 0
`define AXI_HAS_REGIONS_S9 0
`define AXI_HAS_REGIONS_S10 0
`define AXI_HAS_REGIONS_S11 0
`define AXI_HAS_REGIONS_S12 0
`define AXI_HAS_REGIONS_S13 0
`define AXI_HAS_REGIONS_S14 0
`define AXI_HAS_REGIONS_S15 0
`define AXI_HAS_REGIONS_S16 0
`define AXI_HAS_REGIONS 0
`define AXI_BCM_TST_MODE 0
`define AXI_BCM_CDC_INIT 0
`define DWC_NO_TST_MODE
`define DWC_NO_CDC_INIT
`define __GUARD__DW_AXI_CONSTANTS__VH__
`define AXI_BSW 3
`define AXI_BTW 2
`define AXI_LTW ((`AXI_INTERFACE_TYPE >0)? 1 :2)
`define AXI_CTW 4
`define AXI_PTW 3
`define AXI_BRW 2
`define AXI_RRW 2
`define AXI_SW        (`AXI_DW/8)
`define AXI_MAX_NUM_MST_SLVS 17
`define AXI_MAX_NUM_USR_MSTS 16
`define AXI_MAX_NUM_USR_SLVS 16
`define AXI_LT_NORM  2'b00
`define AXI_LT_EX    2'b01
`define AXI_LT_LOCK  2'b10
`define AXI_PT_PRVLGD    3'bxx1
`define AXI_PT_NORM      3'bxx0
`define AXI_PT_SECURE    3'bx1x
`define AXI_PT_NSECURE   3'bx0x
`define AXI_PT_INSTRUCT  3'b1xx
`define AXI_PT_DATA      3'b0xx
`define AXI_PT_PRVLGD_BIT   0
`define AXI_PT_INSTRUCT_BIT 2
`define AXI_RESP_OKAY     2'b00
`define AXI_RESP_EXOKAY   2'b01
`define AXI_RESP_SLVERR   2'b10
`define AXI_RESP_DECERR   2'b11
`define AXI_TMO_COMB  2'b00
`define AXI_TMO_FRWD  2'b01
`define AXI_TMO_FULL  2'b10
`define AXI_NOREQ_LOCKING  0 // No locking functionality required.
`define AXI_REQ_LOCKING    1 // Locking functionality required.
`define AXI_ARB_TYPE_DP   0
`define AXI_ARB_TYPE_FCFS 1
`define AXI_ARB_TYPE_2T   2
`define AXI_ARB_TYPE_USER 3
`define AXI_ARB_TYPE_QOS  4
`define AXI_W_CH 1      // This channel is a write data channel.
`define AXI_NOT_W_CH  0 // This channel is not a write data channel.
`define AXI_AW_CH 1      // This channel is a write address channel.
`define AXI_NOT_AW_CH  0 // This channel is not a write address channel.
`define AXI_R_CH 1      // This channel is a read data channel.
`define AXI_NOT_R_CH  0 // This channel is not a read data channel.
`define AXI_ADDR_CH 1     // This channel is an address channel.
`define AXI_NOT_ADDR_CH 0 // This channel is not an address channel.
`define USE_INT_GI  1 // Use internal grant index.
`define USE_EXT_GI  0 // Use external grant index.
`define AXI_SHARED 1
`define AXI_NOT_SHARED 0
`define AXI_HOLD_VLD_OTHER_S_W (`AXI_NUM_MASTERS*(`AXI_NSP1-1))
`define AXI_HOLD_VLD_OTHER_M_W ((`AXI_NUM_MASTERS > 1) ? (`AXI_NSP1*(`AXI_NUM_MASTERS-1)) : 1)
`define AXI_ARPYLD_PROT_RHS 0
`define AXI_ARPYLD_PROT_LHS ((`AXI_PTW-1) + `AXI_ARPYLD_PROT_RHS)
`define AXI_ARPYLD_PROT    1 
`define AXI_ARPYLD_CACHE_RHS (`AXI_ARPYLD_PROT_LHS + 1)
`define AXI_ARPYLD_CACHE_LHS ((`AXI_CTW-1) + `AXI_ARPYLD_CACHE_RHS)
`define AXI_ARPYLD_CACHE     `AXI_ARPYLD_CACHE_LHS:`AXI_ARPYLD_CACHE_RHS
`define AXI_ARPYLD_LOCK_RHS (`AXI_ARPYLD_CACHE_LHS + 1)
`define AXI_ARPYLD_LOCK_LHS ((`AXI_LTW-1) + `AXI_ARPYLD_LOCK_RHS)
`define AXI_ARPYLD_LOCK     `AXI_ARPYLD_LOCK_LHS:`AXI_ARPYLD_LOCK_RHS
`define AXI_ARPYLD_BURST_RHS (`AXI_ARPYLD_LOCK_LHS + 1)
`define AXI_ARPYLD_BURST_LHS ((`AXI_BTW-1) + `AXI_ARPYLD_BURST_RHS)
`define AXI_ARPYLD_BURST     `AXI_ARPYLD_BURST_LHS:`AXI_ARPYLD_BURST_RHS
`define AXI_ARPYLD_SIZE_RHS (`AXI_ARPYLD_BURST_LHS + 1)
`define AXI_ARPYLD_SIZE_LHS ((`AXI_BSW-1) + `AXI_ARPYLD_SIZE_RHS)
`define AXI_ARPYLD_SIZE     `AXI_ARPYLD_SIZE_LHS:`AXI_ARPYLD_SIZE_RHS
`define AXI_ARPYLD_LEN_RHS (`AXI_ARPYLD_SIZE_LHS + 1)
`define AXI_ARPYLD_LEN_LHS ((`AXI_BLW-1) + `AXI_ARPYLD_LEN_RHS)
`define AXI_ARPYLD_LEN     `AXI_ARPYLD_LEN_LHS:`AXI_ARPYLD_LEN_RHS
`define AXI_ARPYLD_ADDR_RHS (`AXI_ARPYLD_LEN_LHS + 1)
`define AXI_ARPYLD_ADDR_LHS ((`AXI_AW-1) + `AXI_ARPYLD_ADDR_RHS)
`define AXI_ARPYLD_ADDR     `AXI_ARPYLD_ADDR_LHS:`AXI_ARPYLD_ADDR_RHS
`define AXI_ARPYLD_ID_RHS_M (`AXI_ARPYLD_ADDR_LHS + 1)
`define AXI_ARPYLD_ID_LHS_M ((`AXI_MIDW-1) + `AXI_ARPYLD_ID_RHS_M)
`define AXI_ARPYLD_ID_M     `AXI_ARPYLD_ID_LHS_M:`AXI_ARPYLD_ID_RHS_M
`define AXI_ARPYLD_ID_RHS_S (`AXI_ARPYLD_ADDR_LHS + 1)
`define AXI_ARPYLD_ID_LHS_S ((`AXI_SIDW-1) + `AXI_ARPYLD_ID_RHS_S)
`define AXI_ARPYLD_ID_S     `AXI_ARPYLD_ID_LHS_S:`AXI_ARPYLD_ID_RHS_S
`define AXI_RPYLD_LAST_LHS 0
`define AXI_RPYLD_LAST     `AXI_RPYLD_LAST_LHS
`define AXI_RPYLD_RESP_RHS (`AXI_RPYLD_LAST_LHS + 1)
`define AXI_RPYLD_RESP_LHS ((`AXI_RRW-1) + `AXI_RPYLD_RESP_RHS)
`define AXI_RPYLD_RESP     `AXI_RPYLD_RESP_LHS:`AXI_RPYLD_RESP_RHS
`define AXI_RPYLD_DATA_RHS (`AXI_RPYLD_RESP_LHS + 1)
`define AXI_RPYLD_DATA_LHS ((`AXI_DW-1) + `AXI_RPYLD_DATA_RHS)
`define AXI_RPYLD_DATA     `AXI_RPYLD_DATA_LHS:`AXI_RPYLD_DATA_RHS
`define AXI_RPYLD_ID_RHS_M (`AXI_RPYLD_DATA_LHS + 1)
`define AXI_RPYLD_ID_LHS_M ((`AXI_MIDW-1) + `AXI_RPYLD_ID_RHS_M)
`define AXI_RPYLD_ID_M     `AXI_RPYLD_ID_LHS_M:`AXI_RPYLD_ID_RHS_M
`define AXI_RPYLD_ID_RHS_S (`AXI_RPYLD_DATA_LHS + 1)
`define AXI_RPYLD_ID_LHS_S ((`AXI_SIDW-1) + `AXI_RPYLD_ID_RHS_S)
`define AXI_RPYLD_ID_S     `AXI_RPYLD_ID_LHS_S:`AXI_RPYLD_ID_RHS_S
`define AXI_AWPYLD_PROT_RHS 0
`define AXI_AWPYLD_PROT_LHS ((`AXI_PTW-1) + `AXI_AWPYLD_PROT_RHS)
`define AXI_AWPYLD_PROT     `AXI_AWPYLD_PROT_LHS:`AXI_AWPYLD_PROT_RHS
`define AXI_AWPYLD_CACHE_RHS (`AXI_AWPYLD_PROT_LHS + 1)
`define AXI_AWPYLD_CACHE_LHS ((`AXI_CTW-1) + `AXI_AWPYLD_CACHE_RHS)
`define AXI_AWPYLD_CACHE     `AXI_AWPYLD_CACHE_LHS:`AXI_AWPYLD_CACHE_RHS
`define AXI_AWPYLD_LOCK_RHS (`AXI_AWPYLD_CACHE_LHS + 1)
`define AXI_AWPYLD_LOCK_LHS ((`AXI_LTW-1) + `AXI_AWPYLD_LOCK_RHS)
`define AXI_AWPYLD_LOCK     `AXI_AWPYLD_LOCK_LHS:`AXI_AWPYLD_LOCK_RHS
`define AXI_AWPYLD_BURST_RHS (`AXI_AWPYLD_LOCK_LHS + 1)
`define AXI_AWPYLD_BURST_LHS ((`AXI_BTW-1) + `AXI_AWPYLD_BURST_RHS)
`define AXI_AWPYLD_BURST     `AXI_AWPYLD_BURST_LHS:`AXI_AWPYLD_BURST_RHS
`define AXI_AWPYLD_SIZE_RHS (`AXI_AWPYLD_BURST_LHS + 1)
`define AXI_AWPYLD_SIZE_LHS ((`AXI_BSW-1) + `AXI_AWPYLD_SIZE_RHS)
`define AXI_AWPYLD_SIZE     `AXI_AWPYLD_SIZE_LHS:`AXI_AWPYLD_SIZE_RHS
`define AXI_AWPYLD_LEN_RHS (`AXI_AWPYLD_SIZE_LHS + 1)
`define AXI_AWPYLD_LEN_LHS ((`AXI_BLW-1) + `AXI_AWPYLD_LEN_RHS)
`define AXI_AWPYLD_LEN     `AXI_AWPYLD_LEN_LHS:`AXI_AWPYLD_LEN_RHS
`define AXI_AWPYLD_ADDR_RHS (`AXI_AWPYLD_LEN_LHS + 1)
`define AXI_AWPYLD_ADDR_LHS ((`AXI_AW-1) + `AXI_AWPYLD_ADDR_RHS)
`define AXI_AWPYLD_ADDR     `AXI_AWPYLD_ADDR_LHS:`AXI_AWPYLD_ADDR_RHS
`define AXI_AWPYLD_ID_RHS_M (`AXI_AWPYLD_ADDR_LHS + 1)
`define AXI_AWPYLD_ID_LHS_M ((`AXI_MIDW-1) + `AXI_AWPYLD_ID_RHS_M)
`define AXI_AWPYLD_ID_M     `AXI_AWPYLD_ID_LHS_M:`AXI_AWPYLD_ID_RHS_M
`define AXI_AWPYLD_ID_RHS_S (`AXI_AWPYLD_ADDR_LHS + 1)
`define AXI_AWPYLD_ID_LHS_S ((`AXI_SIDW-1) + `AXI_AWPYLD_ID_RHS_S)
`define AXI_AWPYLD_ID_S     `AXI_AWPYLD_ID_LHS_S:`AXI_AWPYLD_ID_RHS_S
`define AXI_WPYLD_LAST_LHS 0
`define AXI_WPYLD_LAST     `AXI_WPYLD_LAST_LHS
`define AXI_WPYLD_STRB_RHS (`AXI_WPYLD_LAST_LHS + 1)
`define AXI_WPYLD_STRB_LHS ((`AXI_SW-1) + `AXI_WPYLD_STRB_RHS)
`define AXI_WPYLD_STRB     `AXI_WPYLD_STRB_LHS:`AXI_WPYLD_STRB_RHS
`define AXI_WPYLD_DATA_RHS (`AXI_WPYLD_STRB_LHS + 1)
`define AXI_WPYLD_DATA_LHS ((`AXI_DW-1) + `AXI_WPYLD_DATA_RHS)
`define AXI_WPYLD_DATA     `AXI_WPYLD_DATA_LHS:`AXI_WPYLD_DATA_RHS
`define AXI_WPYLD_ID_RHS_M (`AXI_WPYLD_DATA_LHS + 1)
`define AXI_WPYLD_ID_LHS_M ((`AXI_MIDW-1) + `AXI_WPYLD_ID_RHS_M)
`define AXI_WPYLD_ID_M     `AXI_WPYLD_ID_LHS_M:`AXI_WPYLD_ID_RHS_M
`define AXI_WPYLD_ID_RHS_S (`AXI_WPYLD_DATA_LHS + 1)
`define AXI_WPYLD_ID_LHS_S ((`AXI_SIDW-1) + `AXI_WPYLD_ID_RHS_S)
`define AXI_WPYLD_ID_S     `AXI_WPYLD_ID_LHS_S:`AXI_WPYLD_ID_RHS_S
`define AXI_BPYLD_RESP_RHS 0
`define AXI_BPYLD_RESP_LHS ((`AXI_BRW-1) + `AXI_BPYLD_RESP_RHS)
`define AXI_BPYLD_RESP     `AXI_BPYLD_RESP_LHS:`AXI_BPYLD_RESP_RHS
`define AXI_BPYLD_ID_RHS_M (`AXI_BPYLD_RESP_LHS + 1)
`define AXI_BPYLD_ID_LHS_M ((`AXI_MIDW-1) + `AXI_BPYLD_ID_RHS_M)
`define AXI_BPYLD_ID_M     `AXI_BPYLD_ID_LHS_M:`AXI_BPYLD_ID_RHS_M
`define AXI_BPYLD_ID_RHS_S (`AXI_BPYLD_RESP_LHS + 1)
`define AXI_BPYLD_ID_LHS_S ((`AXI_SIDW-1) + `AXI_BPYLD_ID_RHS_S)
`define AXI_BPYLD_ID_S     `AXI_BPYLD_ID_LHS_S:`AXI_BPYLD_ID_RHS_S
`define AXI_QOSW  4
`define IC_ADDR_SLICE_LHS  5
`define MAX_APB_DATA_WIDTH 32
`define REG_XCT_RATE_W      12
`define REG_BURSTINESS_W    8
`define REG_PEAK_RATE_W     12
`define APB_ADDR_WIDTH      32
`define AXI_ALSW 4 
`define AXI_ALDW 2
`define AXI_ALBW 2
`define AXI_REGIONW 4
`define PL_BUF_AW 0
`define PL_BUF_AR 0
`define ACT_ID_BUF_POINTER_W_AW_M1 70
`define LOG2_ACT_ID_BUF_POINTER_W_AW_M1 4
`define ACT_ID_BUF_POINTER_W_AR_M1 40
`define LOG2_ACT_ID_BUF_POINTER_W_AR_M1 3
`define ACT_ID_BUF_POINTER_W_AW_M2 70
`define LOG2_ACT_ID_BUF_POINTER_W_AW_M2 4
`define ACT_ID_BUF_POINTER_W_AR_M2 40
`define LOG2_ACT_ID_BUF_POINTER_W_AR_M2 3
`define ACT_ID_BUF_POINTER_W_AW_M3 10
`define LOG2_ACT_ID_BUF_POINTER_W_AW_M3 1
`define ACT_ID_BUF_POINTER_W_AR_M3 40
`define LOG2_ACT_ID_BUF_POINTER_W_AR_M3 3
`define ACT_ID_BUF_POINTER_W_AW_M4 10
`define LOG2_ACT_ID_BUF_POINTER_W_AW_M4 1
`define ACT_ID_BUF_POINTER_W_AR_M4 40
`define LOG2_ACT_ID_BUF_POINTER_W_AR_M4 3
`define ACT_ID_BUF_POINTER_W_AW_M5 10
`define LOG2_ACT_ID_BUF_POINTER_W_AW_M5 1
`define ACT_ID_BUF_POINTER_W_AR_M5 40
`define LOG2_ACT_ID_BUF_POINTER_W_AR_M5 3
`define ACT_ID_BUF_POINTER_W_AW_M6 10
`define LOG2_ACT_ID_BUF_POINTER_W_AW_M6 1
`define ACT_ID_BUF_POINTER_W_AR_M6 40
`define LOG2_ACT_ID_BUF_POINTER_W_AR_M6 3
`define ACT_ID_BUF_POINTER_W_AW_M7 10
`define LOG2_ACT_ID_BUF_POINTER_W_AW_M7 1
`define ACT_ID_BUF_POINTER_W_AR_M7 40
`define LOG2_ACT_ID_BUF_POINTER_W_AR_M7 3
`define ACT_ID_BUF_POINTER_W_AW_M8 10
`define LOG2_ACT_ID_BUF_POINTER_W_AW_M8 1
`define ACT_ID_BUF_POINTER_W_AR_M8 40
`define LOG2_ACT_ID_BUF_POINTER_W_AR_M8 3
`define ACT_ID_BUF_POINTER_W_AW_M9 10
`define LOG2_ACT_ID_BUF_POINTER_W_AW_M9 1
`define ACT_ID_BUF_POINTER_W_AR_M9 40
`define LOG2_ACT_ID_BUF_POINTER_W_AR_M9 3
`define ACT_ID_BUF_POINTER_W_AW_M10 10
`define LOG2_ACT_ID_BUF_POINTER_W_AW_M10 1
`define ACT_ID_BUF_POINTER_W_AR_M10 40
`define LOG2_ACT_ID_BUF_POINTER_W_AR_M10 3
`define ACT_ID_BUF_POINTER_W_AW_M11 10
`define LOG2_ACT_ID_BUF_POINTER_W_AW_M11 1
`define ACT_ID_BUF_POINTER_W_AR_M11 40
`define LOG2_ACT_ID_BUF_POINTER_W_AR_M11 3
`define ACT_ID_BUF_POINTER_W_AW_M12 10
`define LOG2_ACT_ID_BUF_POINTER_W_AW_M12 1
`define ACT_ID_BUF_POINTER_W_AR_M12 40
`define LOG2_ACT_ID_BUF_POINTER_W_AR_M12 3
`define ACT_ID_BUF_POINTER_W_AW_M13 10
`define LOG2_ACT_ID_BUF_POINTER_W_AW_M13 1
`define ACT_ID_BUF_POINTER_W_AR_M13 40
`define LOG2_ACT_ID_BUF_POINTER_W_AR_M13 3
`define ACT_ID_BUF_POINTER_W_AW_M14 10
`define LOG2_ACT_ID_BUF_POINTER_W_AW_M14 1
`define ACT_ID_BUF_POINTER_W_AR_M14 40
`define LOG2_ACT_ID_BUF_POINTER_W_AR_M14 3
`define ACT_ID_BUF_POINTER_W_AW_M15 10
`define LOG2_ACT_ID_BUF_POINTER_W_AW_M15 1
`define ACT_ID_BUF_POINTER_W_AR_M15 40
`define LOG2_ACT_ID_BUF_POINTER_W_AR_M15 3
`define ACT_ID_BUF_POINTER_W_AW_M16 10
`define LOG2_ACT_ID_BUF_POINTER_W_AW_M16 1
`define ACT_ID_BUF_POINTER_W_AR_M16 40
`define LOG2_ACT_ID_BUF_POINTER_W_AR_M16 3
`define AXI_HAS_WID (`AXI_INTERFACE_TYPE==0)
