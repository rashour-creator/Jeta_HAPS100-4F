//##########################################################
// Generated undef unprefix file for workspace: DW_axi_a2x
//##########################################################

`ifdef __GUARD__DW_AXI_A2X_DEFINE_CONSTANTS__VH__
  `undef __GUARD__DW_AXI_A2X_DEFINE_CONSTANTS__VH__
`endif 

`ifdef A2X_BSW
  `undef A2X_BSW
`endif 

`ifdef A2X_BTW
  `undef A2X_BTW
`endif 

`ifdef A2X_LTW
  `undef A2X_LTW
`endif 

`ifdef A2X_CTW
  `undef A2X_CTW
`endif 

`ifdef A2X_PTW
  `undef A2X_PTW
`endif 

`ifdef A2X_RSW
  `undef A2X_RSW
`endif 

`ifdef A2X_BRESPW
  `undef A2X_BRESPW
`endif 

`ifdef A2X_RRESPW
  `undef A2X_RRESPW
`endif 

`ifdef A2X_HIDW
  `undef A2X_HIDW
`endif 

`ifdef A2X_HBLW
  `undef A2X_HBLW
`endif 

`ifdef A2X_HBTYPE_W
  `undef A2X_HBTYPE_W
`endif 

`ifdef A2X_MAX_BSBW
  `undef A2X_MAX_BSBW
`endif 

`ifdef CT_MODE
  `undef CT_MODE
`endif 

`ifdef SNF_MODE
  `undef SNF_MODE
`endif 

`ifdef ABURST_FIXED
  `undef ABURST_FIXED
`endif 

`ifdef ABURST_INCR
  `undef ABURST_INCR
`endif 

`ifdef ABURST_WRAP
  `undef ABURST_WRAP
`endif 

`ifdef HTRANS_IDLE
  `undef HTRANS_IDLE
`endif 

`ifdef HTRANS_BUSY
  `undef HTRANS_BUSY
`endif 

`ifdef HTRANS_NSEQ
  `undef HTRANS_NSEQ
`endif 

`ifdef HTRANS_SEQ
  `undef HTRANS_SEQ
`endif 

`ifdef HBURST_SINGLE
  `undef HBURST_SINGLE
`endif 

`ifdef HBURST_INCR
  `undef HBURST_INCR
`endif 

`ifdef HBURST_WRAP4
  `undef HBURST_WRAP4
`endif 

`ifdef HBURST_INCR4
  `undef HBURST_INCR4
`endif 

`ifdef HBURST_WRAP8
  `undef HBURST_WRAP8
`endif 

`ifdef HBURST_INCR8
  `undef HBURST_INCR8
`endif 

`ifdef HBURST_WRAP16
  `undef HBURST_WRAP16
`endif 

`ifdef HBURST_INCR16
  `undef HBURST_INCR16
`endif 

`ifdef HSIZE_8
  `undef HSIZE_8
`endif 

`ifdef HSIZE_16
  `undef HSIZE_16
`endif 

`ifdef HSIZE_32
  `undef HSIZE_32
`endif 

`ifdef HSIZE_64
  `undef HSIZE_64
`endif 

`ifdef HSIZE_128
  `undef HSIZE_128
`endif 

`ifdef HSIZE_256
  `undef HSIZE_256
`endif 

`ifdef HSIZE_512
  `undef HSIZE_512
`endif 

`ifdef HSIZE_1024
  `undef HSIZE_1024
`endif 

`ifdef HSIZE_8BIT
  `undef HSIZE_8BIT
`endif 

`ifdef HSIZE_16BIT
  `undef HSIZE_16BIT
`endif 

`ifdef HSIZE_32BIT
  `undef HSIZE_32BIT
`endif 

`ifdef HSIZE_64BIT
  `undef HSIZE_64BIT
`endif 

`ifdef HSIZE_128BIT
  `undef HSIZE_128BIT
`endif 

`ifdef HSIZE_256BIT
  `undef HSIZE_256BIT
`endif 

`ifdef HSIZE_512BIT
  `undef HSIZE_512BIT
`endif 

`ifdef HSIZE_1024BIT
  `undef HSIZE_1024BIT
`endif 

`ifdef HSIZE_BYTE
  `undef HSIZE_BYTE
`endif 

`ifdef HSIZE_WORD16
  `undef HSIZE_WORD16
`endif 

`ifdef HSIZE_WORD32
  `undef HSIZE_WORD32
`endif 

`ifdef HSIZE_WORD64
  `undef HSIZE_WORD64
`endif 

`ifdef HSIZE_WORD128
  `undef HSIZE_WORD128
`endif 

`ifdef HSIZE_WORD256
  `undef HSIZE_WORD256
`endif 

`ifdef HSIZE_WORD512
  `undef HSIZE_WORD512
`endif 

`ifdef HSIZE_WORD1024
  `undef HSIZE_WORD1024
`endif 

`ifdef HPROT_DATA
  `undef HPROT_DATA
`endif 

`ifdef HPROT_PRIV
  `undef HPROT_PRIV
`endif 

`ifdef HPROT_BUFF
  `undef HPROT_BUFF
`endif 

`ifdef HPROT_CACHE
  `undef HPROT_CACHE
`endif 

`ifdef HRESP_OKAY
  `undef HRESP_OKAY
`endif 

`ifdef HRESP_ERROR
  `undef HRESP_ERROR
`endif 

`ifdef HRESP_RETRY
  `undef HRESP_RETRY
`endif 

`ifdef HRESP_SPLIT
  `undef HRESP_SPLIT
`endif 

`ifdef AFIXED
  `undef AFIXED
`endif 

`ifdef AINCR
  `undef AINCR
`endif 

`ifdef AWRAP
  `undef AWRAP
`endif 

`ifdef AOKAY
  `undef AOKAY
`endif 

`ifdef AEXOKAY
  `undef AEXOKAY
`endif 

`ifdef ASLVERR
  `undef ASLVERR
`endif 

`ifdef ADECERR
  `undef ADECERR
`endif 

`ifdef __GUARD__DW_AXI_A2X_CC_CONSTANTS__VH__
  `undef __GUARD__DW_AXI_A2X_CC_CONSTANTS__VH__
`endif 

`ifdef USE_FOUNDATION
  `undef USE_FOUNDATION
`endif 

`ifdef A2X_USE_FOUNDATION
  `undef A2X_USE_FOUNDATION
`endif 

`ifdef A2X_LOWPWR_IF
  `undef A2X_LOWPWR_IF
`endif 

`ifdef A2X_LOWPWR_NOPX_CNT
  `undef A2X_LOWPWR_NOPX_CNT
`endif 

`ifdef A2X_PP_MODE
  `undef A2X_PP_MODE
`endif 

`ifdef A2X_AHB_INTERFACE_TYPE
  `undef A2X_AHB_INTERFACE_TYPE
`endif 

`ifdef A2X_HAS_EXTD_MEMTYPE
  `undef A2X_HAS_EXTD_MEMTYPE
`endif 

`ifdef A2X_HAS_SECURE_XFER
  `undef A2X_HAS_SECURE_XFER
`endif 

`ifdef A2X_HAS_EXCL_XFER
  `undef A2X_HAS_EXCL_XFER
`endif 

`ifdef A2X_HPTW
  `undef A2X_HPTW
`endif 

`ifdef A2X_AXI_INTERFACE_TYPE
  `undef A2X_AXI_INTERFACE_TYPE
`endif 

`ifdef A2X_INT_AXI3
  `undef A2X_INT_AXI3
`endif 

`ifdef A2X_INT_LTW
  `undef A2X_INT_LTW
`endif 

`ifdef A2X_HAS_AXI3
  `undef A2X_HAS_AXI3
`endif 

`ifdef A2X_HAS_AXI4
  `undef A2X_HAS_AXI4
`endif 

`ifdef A2X_HAS_ACELITE
  `undef A2X_HAS_ACELITE
`endif 

`ifdef A2X_AHB_LITE_MODE
  `undef A2X_AHB_LITE_MODE
`endif 

`ifdef A2X_AHB_SCALAR_HRESP
  `undef A2X_AHB_SCALAR_HRESP
`endif 

`ifdef A2X_AHB_SPLIT_MODE
  `undef A2X_AHB_SPLIT_MODE
`endif 

`ifdef AHB_SPLIT_MODE
  `undef AHB_SPLIT_MODE
`endif 

`ifdef A2X_NUM_AHBM
  `undef A2X_NUM_AHBM
`endif 

`ifdef A2X_HREADY_LOW_PERIOD
  `undef A2X_HREADY_LOW_PERIOD
`endif 

`ifdef A2X_LOCKED
  `undef A2X_LOCKED
`endif 

`ifdef A2X_CLK_MODE
  `undef A2X_CLK_MODE
`endif 

`ifdef A2X_PP_SYNC_DEPTH
  `undef A2X_PP_SYNC_DEPTH
`endif 

`ifdef F_SYNC_TYPE_PP
  `undef F_SYNC_TYPE_PP
`endif 

`ifdef A2X_SP_SYNC_DEPTH
  `undef A2X_SP_SYNC_DEPTH
`endif 

`ifdef F_SYNC_TYPE_SP
  `undef F_SYNC_TYPE_SP
`endif 

`ifdef A2X_SYNC_DEPTH_BUSY
  `undef A2X_SYNC_DEPTH_BUSY
`endif 

`ifdef A2X_PP_IDW
  `undef A2X_PP_IDW
`endif 

`ifdef A2X_IDW
  `undef A2X_IDW
`endif 

`ifdef A2X_SP_IDW
  `undef A2X_SP_IDW
`endif 

`ifdef A2X_PP_AW
  `undef A2X_PP_AW
`endif 

`ifdef A2X_AW
  `undef A2X_AW
`endif 

`ifdef A2X_SP_AW
  `undef A2X_SP_AW
`endif 

`ifdef A2X_BOUNDARY_W
  `undef A2X_BOUNDARY_W
`endif 

`ifdef A2X_PP_BLW
  `undef A2X_PP_BLW
`endif 

`ifdef A2X_SP_BLW
  `undef A2X_SP_BLW
`endif 

`ifdef A2X_BLW
  `undef A2X_BLW
`endif 

`ifdef A2X_MAX_ALEN
  `undef A2X_MAX_ALEN
`endif 

`ifdef A2X_PP_DW
  `undef A2X_PP_DW
`endif 

`ifdef A2X_SP_DW
  `undef A2X_SP_DW
`endif 

`ifdef A2X_RS_RATIO
  `undef A2X_RS_RATIO
`endif 

`ifdef A2X_RS_RATIO_LOG2
  `undef A2X_RS_RATIO_LOG2
`endif 

`ifdef A2X_PP_ENDIAN
  `undef A2X_PP_ENDIAN
`endif 

`ifdef A2X_SP_ENDIAN
  `undef A2X_SP_ENDIAN
`endif 

`ifdef A2X_WBUF_MODE
  `undef A2X_WBUF_MODE
`endif 

`ifdef A2X_HCBUF_MODE
  `undef A2X_HCBUF_MODE
`endif 

`ifdef A2X_APB_MODE
  `undef A2X_APB_MODE
`endif 

`ifdef A2X_HCSNF_WLEN
  `undef A2X_HCSNF_WLEN
`endif 

`ifdef A2X_SNF_AWLEN_DFLT
  `undef A2X_SNF_AWLEN_DFLT
`endif 

`ifdef A2X_SNF_AWLEN_MIN
  `undef A2X_SNF_AWLEN_MIN
`endif 

`ifdef A2X_HINCR_HCBCNT
  `undef A2X_HINCR_HCBCNT
`endif 

`ifdef A2X_SINGLE_RBCNT
  `undef A2X_SINGLE_RBCNT
`endif 

`ifdef A2X_SINGLE_WBCNT
  `undef A2X_SINGLE_WBCNT
`endif 

`ifdef A2X_HINCR_WBCNT_MIN
  `undef A2X_HINCR_WBCNT_MIN
`endif 

`ifdef A2X_HINCR_WBCNT_MAX
  `undef A2X_HINCR_WBCNT_MAX
`endif 

`ifdef A2X_HINCR_AWLEN_DFLT
  `undef A2X_HINCR_AWLEN_DFLT
`endif 

`ifdef A2X_HINCR_AWLEN_MIN
  `undef A2X_HINCR_AWLEN_MIN
`endif 

`ifdef A2X_BRESP_MODE
  `undef A2X_BRESP_MODE
`endif 

`ifdef A2X_BRESP_ORDER
  `undef A2X_BRESP_ORDER
`endif 

`ifdef A2X_OSW_EN
  `undef A2X_OSW_EN
`endif 

`ifdef A2X_NUM_UWID
  `undef A2X_NUM_UWID
`endif 

`ifdef A2X_SP_OSAW_LIMIT_P1
  `undef A2X_SP_OSAW_LIMIT_P1
`endif 

`ifdef A2X_SP_OSAW_LIMIT
  `undef A2X_SP_OSAW_LIMIT
`endif 

`ifdef A2X_OSAW_LIMIT
  `undef A2X_OSAW_LIMIT
`endif 

`ifdef A2X_PP_OSAW_LIMIT_P1
  `undef A2X_PP_OSAW_LIMIT_P1
`endif 

`ifdef A2X_PP_OSAW_LIMIT
  `undef A2X_PP_OSAW_LIMIT
`endif 

`ifdef A2X_B_OSW_LIMIT_P1
  `undef A2X_B_OSW_LIMIT_P1
`endif 

`ifdef A2X_B_OSW_LIMIT
  `undef A2X_B_OSW_LIMIT
`endif 

`ifdef A2X_OSW_LIMIT
  `undef A2X_OSW_LIMIT
`endif 

`ifdef A2X_RBUF_MODE
  `undef A2X_RBUF_MODE
`endif 

`ifdef A2X_HCSNF_RLEN
  `undef A2X_HCSNF_RLEN
`endif 

`ifdef A2X_SNF_ARLEN_DFLT
  `undef A2X_SNF_ARLEN_DFLT
`endif 

`ifdef A2X_SNF_ARLEN_MIN
  `undef A2X_SNF_ARLEN_MIN
`endif 

`ifdef A2X_AHB_RRECALL_DEPTH
  `undef A2X_AHB_RRECALL_DEPTH
`endif 

`ifdef A2X_AHB_EBT_MODE
  `undef A2X_AHB_EBT_MODE
`endif 

`ifdef A2X_HINCR_RBCNT_MIN
  `undef A2X_HINCR_RBCNT_MIN
`endif 

`ifdef A2X_HINCR_RBCNT_MAX
  `undef A2X_HINCR_RBCNT_MAX
`endif 

`ifdef A2X_LKMODE_MAX_PREFETCH
  `undef A2X_LKMODE_MAX_PREFETCH
`endif 

`ifdef A2X_HINCR_ARLEN_DFLT
  `undef A2X_HINCR_ARLEN_DFLT
`endif 

`ifdef A2X_HINCR_ARLEN_MIN
  `undef A2X_HINCR_ARLEN_MIN
`endif 

`ifdef A2X_READ_INTLEV
  `undef A2X_READ_INTLEV
`endif 

`ifdef A2X_READ_ORDER
  `undef A2X_READ_ORDER
`endif 

`ifdef SIM_REORDER
  `undef SIM_REORDER
`endif 

`ifdef A2X_OSR_EN
  `undef A2X_OSR_EN
`endif 

`ifdef A2X_NUM_URID
  `undef A2X_NUM_URID
`endif 

`ifdef A2X_OSR_LIMIT_P1
  `undef A2X_OSR_LIMIT_P1
`endif 

`ifdef A2X_OSR_LIMIT
  `undef A2X_OSR_LIMIT
`endif 

`ifdef A2X_A_UBW
  `undef A2X_A_UBW
`endif 

`ifdef A2X_USER_SIGNAL_XFER_MODE
  `undef A2X_USER_SIGNAL_XFER_MODE
`endif 

`ifdef A2X_WUSER_BITS_PER_BYTE
  `undef A2X_WUSER_BITS_PER_BYTE
`endif 

`ifdef A2X_RUSER_BITS_PER_BYTE
  `undef A2X_RUSER_BITS_PER_BYTE
`endif 

`ifdef A2X_W_UBW
  `undef A2X_W_UBW
`endif 

`ifdef A2X_R_UBW
  `undef A2X_R_UBW
`endif 

`ifdef A2X_AWSBW
  `undef A2X_AWSBW
`endif 

`ifdef A2X_ARSBW
  `undef A2X_ARSBW
`endif 

`ifdef A2X_WSBW
  `undef A2X_WSBW
`endif 

`ifdef A2X_RSBW
  `undef A2X_RSBW
`endif 

`ifdef A2X_BSBW
  `undef A2X_BSBW
`endif 

`ifdef A2X_INC_QOS
  `undef A2X_INC_QOS
`endif 

`ifdef A2X_HAS_QOS
  `undef A2X_HAS_QOS
`endif 

`ifdef A2X_INC_REGION
  `undef A2X_INC_REGION
`endif 

`ifdef A2X_HAS_REGION
  `undef A2X_HAS_REGION
`endif 

`ifdef A2X_AW_FIFO_DEPTH
  `undef A2X_AW_FIFO_DEPTH
`endif 

`ifdef A2X_WD_FIFO_DEPTH
  `undef A2X_WD_FIFO_DEPTH
`endif 

`ifdef A2X_BRESP_FIFO_DEPTH
  `undef A2X_BRESP_FIFO_DEPTH
`endif 

`ifdef A2X_AR_FIFO_DEPTH
  `undef A2X_AR_FIFO_DEPTH
`endif 

`ifdef A2X_RD_FIFO_DEPTH
  `undef A2X_RD_FIFO_DEPTH
`endif 

`ifdef A2X_LK_RD_FIFO_DEPTH
  `undef A2X_LK_RD_FIFO_DEPTH
`endif 

`ifdef A2X_AUTO_LINK_SPLIT_MODE
  `undef A2X_AUTO_LINK_SPLIT_MODE
`endif 

`ifdef A2X_AR_SP_PIPELINE
  `undef A2X_AR_SP_PIPELINE
`endif 

`ifdef A2X_AW_SP_PIPELINE
  `undef A2X_AW_SP_PIPELINE
`endif 

`ifdef A2X_RS_AR_TMO
  `undef A2X_RS_AR_TMO
`endif 

`ifdef A2X_RS_AW_TMO
  `undef A2X_RS_AW_TMO
`endif 

`ifdef A2X_RS_R_TMO
  `undef A2X_RS_R_TMO
`endif 

`ifdef A2X_RS_W_TMO
  `undef A2X_RS_W_TMO
`endif 

`ifdef A2X_RS_B_TMO
  `undef A2X_RS_B_TMO
`endif 

`ifdef A2X_AHB_LOCKED
  `undef A2X_AHB_LOCKED
`endif 

`ifdef A2X_HAS_LOCKED
  `undef A2X_HAS_LOCKED
`endif 

`ifdef A2X_INT_NUM_AHBM
  `undef A2X_INT_NUM_AHBM
`endif 

`ifdef A2X_UPSIZE
  `undef A2X_UPSIZE
`endif 

`ifdef A2X_DOWNSIZE
  `undef A2X_DOWNSIZE
`endif 

`ifdef A2X_IS_UPSIZED
  `undef A2X_IS_UPSIZED
`endif 

`ifdef A2X_IS_DOWNSIZED
  `undef A2X_IS_DOWNSIZED
`endif 

`ifdef A2X_HAS_RBUF
  `undef A2X_HAS_RBUF
`endif 

`ifdef A2X_IS_EQSIZED
  `undef A2X_IS_EQSIZED
`endif 

`ifdef A2X_HAS_NBUF_MODE
  `undef A2X_HAS_NBUF_MODE
`endif 

`ifdef A2X_HAS_HINCR_HCBCNT
  `undef A2X_HAS_HINCR_HCBCNT
`endif 

`ifdef A2X_HAS_SINGLE_RBCNT
  `undef A2X_HAS_SINGLE_RBCNT
`endif 

`ifdef A2X_HAS_SINGLE_WBCNT
  `undef A2X_HAS_SINGLE_WBCNT
`endif 

`ifdef A2X_HAS_CNT_M1
  `undef A2X_HAS_CNT_M1
`endif 

`ifdef A2X_HAS_CNT_M2
  `undef A2X_HAS_CNT_M2
`endif 

`ifdef A2X_HAS_CNT_M3
  `undef A2X_HAS_CNT_M3
`endif 

`ifdef A2X_HAS_CNT_M4
  `undef A2X_HAS_CNT_M4
`endif 

`ifdef A2X_HAS_CNT_M5
  `undef A2X_HAS_CNT_M5
`endif 

`ifdef A2X_HAS_CNT_M6
  `undef A2X_HAS_CNT_M6
`endif 

`ifdef A2X_HAS_CNT_M7
  `undef A2X_HAS_CNT_M7
`endif 

`ifdef A2X_HAS_CNT_M8
  `undef A2X_HAS_CNT_M8
`endif 

`ifdef A2X_HAS_CNT_M9
  `undef A2X_HAS_CNT_M9
`endif 

`ifdef A2X_HAS_CNT_M10
  `undef A2X_HAS_CNT_M10
`endif 

`ifdef A2X_HAS_CNT_M11
  `undef A2X_HAS_CNT_M11
`endif 

`ifdef A2X_HAS_CNT_M12
  `undef A2X_HAS_CNT_M12
`endif 

`ifdef A2X_HAS_CNT_M13
  `undef A2X_HAS_CNT_M13
`endif 

`ifdef A2X_HAS_CNT_M14
  `undef A2X_HAS_CNT_M14
`endif 

`ifdef A2X_HAS_CNT_M15
  `undef A2X_HAS_CNT_M15
`endif 

`ifdef A2X_HAS_LOWPWR_IF
  `undef A2X_HAS_LOWPWR_IF
`endif 

`ifdef A2X_HAS_USER_SIGNAL_XFER_MODE
  `undef A2X_HAS_USER_SIGNAL_XFER_MODE
`endif 

`ifdef A2X_INT_HASBW
  `undef A2X_INT_HASBW
`endif 

`ifdef A2X_HAS_HASB
  `undef A2X_HAS_HASB
`endif 

`ifdef A2X_INT_HWSBW
  `undef A2X_INT_HWSBW
`endif 

`ifdef A2X_HAS_HWSB
  `undef A2X_HAS_HWSB
`endif 

`ifdef A2X_INT_HRSBW
  `undef A2X_INT_HRSBW
`endif 

`ifdef A2X_HAS_HRSB
  `undef A2X_HAS_HRSB
`endif 

`ifdef A2X_HAS_AWSB
  `undef A2X_HAS_AWSB
`endif 

`ifdef A2X_INT_AWSBW
  `undef A2X_INT_AWSBW
`endif 

`ifdef A2X_HAS_WSB
  `undef A2X_HAS_WSB
`endif 

`ifdef A2X_INT_WSBW
  `undef A2X_INT_WSBW
`endif 

`ifdef A2X_HAS_ARSB
  `undef A2X_HAS_ARSB
`endif 

`ifdef A2X_INT_ARSBW
  `undef A2X_INT_ARSBW
`endif 

`ifdef A2X_HAS_RSB
  `undef A2X_HAS_RSB
`endif 

`ifdef A2X_INT_RSBW
  `undef A2X_INT_RSBW
`endif 

`ifdef A2X_HAS_BSB
  `undef A2X_HAS_BSB
`endif 

`ifdef A2X_INT_BSBW
  `undef A2X_INT_BSBW
`endif 

`ifdef A2X_PP_IS_AHB
  `undef A2X_PP_IS_AHB
`endif 

`ifdef A2X_PP_IS_AXI
  `undef A2X_PP_IS_AXI
`endif 

`ifdef A2X_CLK_IS_SYNC
  `undef A2X_CLK_IS_SYNC
`endif 

`ifdef A2X_AW_FIFO_DEPTH_LOG2
  `undef A2X_AW_FIFO_DEPTH_LOG2
`endif 

`ifdef A2X_AR_FIFO_DEPTH_LOG2
  `undef A2X_AR_FIFO_DEPTH_LOG2
`endif 

`ifdef A2X_BRESP_FIFO_DEPTH_LOG2
  `undef A2X_BRESP_FIFO_DEPTH_LOG2
`endif 

`ifdef A2X_WD_FIFO_DEPTH_LOG2
  `undef A2X_WD_FIFO_DEPTH_LOG2
`endif 

`ifdef A2X_RD_FIFO_DEPTH_LOG2
  `undef A2X_RD_FIFO_DEPTH_LOG2
`endif 

`ifdef A2X_B_OSW_LIMIT_LOG2
  `undef A2X_B_OSW_LIMIT_LOG2
`endif 

`ifdef A2X_PP_OSAW_LIMIT_LOG2
  `undef A2X_PP_OSAW_LIMIT_LOG2
`endif 

`ifdef A2X_SP_OSAW_LIMIT_LOG2
  `undef A2X_SP_OSAW_LIMIT_LOG2
`endif 

`ifdef A2X_OSR_LIMIT_LOG2
  `undef A2X_OSR_LIMIT_LOG2
`endif 

`ifdef A2X_LK_RD_FIFO_DEPTH_LOG2
  `undef A2X_LK_RD_FIFO_DEPTH_LOG2
`endif 

`ifdef A2X_PP_DW_LOG2
  `undef A2X_PP_DW_LOG2
`endif 

`ifdef A2X_SP_DW_LOG2
  `undef A2X_SP_DW_LOG2
`endif 

`ifdef A2X_PP_NUM_BYTES
  `undef A2X_PP_NUM_BYTES
`endif 

`ifdef A2X_PP_WSTRB_DW
  `undef A2X_PP_WSTRB_DW
`endif 

`ifdef A2X_SP_NUM_BYTES
  `undef A2X_SP_NUM_BYTES
`endif 

`ifdef A2X_SP_WSTRB_DW
  `undef A2X_SP_WSTRB_DW
`endif 

`ifdef A2X_PP_MAX_SIZE
  `undef A2X_PP_MAX_SIZE
`endif 

`ifdef A2X_SP_MAX_SIZE
  `undef A2X_SP_MAX_SIZE
`endif 

`ifdef A2X_MAX_PP_TOTAL_BYTES
  `undef A2X_MAX_PP_TOTAL_BYTES
`endif 

`ifdef A2X_MAX_SP_TOTAL_BYTES
  `undef A2X_MAX_SP_TOTAL_BYTES
`endif 

`ifdef A2X_MAX_TOTAL_BYTES
  `undef A2X_MAX_TOTAL_BYTES
`endif 

`ifdef A2X_MAX_TOTAL_BYTES_LOG2
  `undef A2X_MAX_TOTAL_BYTES_LOG2
`endif 

`ifdef A2X_PP_NUM_BYTES_LOG2
  `undef A2X_PP_NUM_BYTES_LOG2
`endif 

`ifdef A2X_SP_NUM_BYTES_LOG2
  `undef A2X_SP_NUM_BYTES_LOG2
`endif 

`ifdef A2X_PP_DW_16
  `undef A2X_PP_DW_16
`endif 

`ifdef A2X_PP_DW_32
  `undef A2X_PP_DW_32
`endif 

`ifdef A2X_PP_DW_64
  `undef A2X_PP_DW_64
`endif 

`ifdef A2X_PP_DW_128
  `undef A2X_PP_DW_128
`endif 

`ifdef A2X_PP_DW_256
  `undef A2X_PP_DW_256
`endif 

`ifdef A2X_PP_DW_512
  `undef A2X_PP_DW_512
`endif 

`ifdef A2X_PP_DW_1024
  `undef A2X_PP_DW_1024
`endif 

`ifdef A2X_SP_DW_32
  `undef A2X_SP_DW_32
`endif 

`ifdef A2X_SP_DW_64
  `undef A2X_SP_DW_64
`endif 

`ifdef A2X_SP_DW_128
  `undef A2X_SP_DW_128
`endif 

`ifdef A2X_SP_DW_256
  `undef A2X_SP_DW_256
`endif 

`ifdef A2X_SP_DW_512
  `undef A2X_SP_DW_512
`endif 

`ifdef A2X_SP_DW_1024
  `undef A2X_SP_DW_1024
`endif 

`ifdef A2X_DS_RATIO_2
  `undef A2X_DS_RATIO_2
`endif 

`ifdef A2X_DS_RATIO_4
  `undef A2X_DS_RATIO_4
`endif 

`ifdef A2X_DS_RATIO_8
  `undef A2X_DS_RATIO_8
`endif 

`ifdef DWC_NO_TST_MODE
  `undef DWC_NO_TST_MODE
`endif 

`ifdef DWC_NO_CDC_INIT
  `undef DWC_NO_CDC_INIT
`endif 

`ifdef A2X_SIM_SEED
  `undef A2X_SIM_SEED
`endif 

`ifdef A2X_SIM_APB_CLK_PERIOD
  `undef A2X_SIM_APB_CLK_PERIOD
`endif 

`ifdef A2X_SIM_PP_CLK_PERIOD
  `undef A2X_SIM_PP_CLK_PERIOD
`endif 

`ifdef A2X_SIM_SP_CLK_PERIOD
  `undef A2X_SIM_SP_CLK_PERIOD
`endif 

`ifdef A2X_SP_CLK_SKEW
  `undef A2X_SP_CLK_SKEW
`endif 

`ifdef A2X_INACTIVE_VAL
  `undef A2X_INACTIVE_VAL
`endif 

`ifdef A2X_ASYNC_CLKS
  `undef A2X_ASYNC_CLKS
`endif 

`ifdef A2X_DUAL_CLK
  `undef A2X_DUAL_CLK
`endif 

`ifdef A2X_N_TESTCASE_DUPLICATION
  `undef A2X_N_TESTCASE_DUPLICATION
`endif 

`ifdef A2X_PRIMEPOWER_SIM
  `undef A2X_PRIMEPOWER_SIM
`endif 

`ifdef A2X_SIM_IS_PRIMEPOWER
  `undef A2X_SIM_IS_PRIMEPOWER
`endif 

`ifdef A2X_VERIF_EN
  `undef A2X_VERIF_EN
`endif 

`ifdef A2X_HRESPW
  `undef A2X_HRESPW
`endif 

`ifdef A2X_HRESP_WIDTH_2
  `undef A2X_HRESP_WIDTH_2
`endif 

`ifdef __GUARD__DW_AXI_A2X_BCM_PARAMS__VH__
  `undef __GUARD__DW_AXI_A2X_BCM_PARAMS__VH__
`endif 

`ifdef DW_AXI_A2X_RM_BCM00_AND
  `undef DW_AXI_A2X_RM_BCM00_AND
`endif 

`ifdef DW_AXI_A2X_RM_BCM00_ATPG_MX
  `undef DW_AXI_A2X_RM_BCM00_ATPG_MX
`endif 

`ifdef DW_AXI_A2X_RM_BCM00_CK_AND
  `undef DW_AXI_A2X_RM_BCM00_CK_AND
`endif 

`ifdef DW_AXI_A2X_RM_BCM00_CK_BUF
  `undef DW_AXI_A2X_RM_BCM00_CK_BUF
`endif 

`ifdef DW_AXI_A2X_RM_BCM00_CK_GT_LAT
  `undef DW_AXI_A2X_RM_BCM00_CK_GT_LAT
`endif 

`ifdef DW_AXI_A2X_RM_BCM00_CK_MX
  `undef DW_AXI_A2X_RM_BCM00_CK_MX
`endif 

`ifdef DW_AXI_A2X_RM_BCM00_CK_OR
  `undef DW_AXI_A2X_RM_BCM00_CK_OR
`endif 

`ifdef DW_AXI_A2X_RM_BCM00_MAJ
  `undef DW_AXI_A2X_RM_BCM00_MAJ
`endif 

`ifdef DW_AXI_A2X_RM_BCM00_MX
  `undef DW_AXI_A2X_RM_BCM00_MX
`endif 

`ifdef DW_AXI_A2X_RM_BCM00_OR
  `undef DW_AXI_A2X_RM_BCM00_OR
`endif 

`ifdef DW_AXI_A2X_RM_BCM01
  `undef DW_AXI_A2X_RM_BCM01
`endif 

`ifdef DW_AXI_A2X_RM_BCM02
  `undef DW_AXI_A2X_RM_BCM02
`endif 

`ifdef DW_AXI_A2X_RM_BCM03
  `undef DW_AXI_A2X_RM_BCM03
`endif 

`ifdef DW_AXI_A2X_RM_BCM04
  `undef DW_AXI_A2X_RM_BCM04
`endif 

`ifdef DW_AXI_A2X_RM_BCM05
  `undef DW_AXI_A2X_RM_BCM05
`endif 

`ifdef DW_AXI_A2X_RM_BCM05_ATV
  `undef DW_AXI_A2X_RM_BCM05_ATV
`endif 

`ifdef DW_AXI_A2X_RM_BCM05_CF
  `undef DW_AXI_A2X_RM_BCM05_CF
`endif 

`ifdef DW_AXI_A2X_RM_BCM05_EF
  `undef DW_AXI_A2X_RM_BCM05_EF
`endif 

`ifdef DW_AXI_A2X_RM_BCM05_EF_ATV
  `undef DW_AXI_A2X_RM_BCM05_EF_ATV
`endif 

`ifdef DW_AXI_A2X_RM_BCM06
  `undef DW_AXI_A2X_RM_BCM06
`endif 

`ifdef DW_AXI_A2X_RM_BCM06_ATV
  `undef DW_AXI_A2X_RM_BCM06_ATV
`endif 

`ifdef DW_AXI_A2X_RM_BCM07
  `undef DW_AXI_A2X_RM_BCM07
`endif 

`ifdef DW_AXI_A2X_RM_BCM07_ATV
  `undef DW_AXI_A2X_RM_BCM07_ATV
`endif 

`ifdef DW_AXI_A2X_RM_BCM07_EF
  `undef DW_AXI_A2X_RM_BCM07_EF
`endif 

`ifdef DW_AXI_A2X_RM_BCM07_EF_ATV
  `undef DW_AXI_A2X_RM_BCM07_EF_ATV
`endif 

`ifdef DW_AXI_A2X_RM_BCM07_EFES
  `undef DW_AXI_A2X_RM_BCM07_EFES
`endif 

`ifdef DW_AXI_A2X_RM_BCM07_RS
  `undef DW_AXI_A2X_RM_BCM07_RS
`endif 

`ifdef DW_AXI_A2X_RM_BCM08
  `undef DW_AXI_A2X_RM_BCM08
`endif 

`ifdef DW_AXI_A2X_RM_BCM09
  `undef DW_AXI_A2X_RM_BCM09
`endif 

`ifdef DW_AXI_A2X_RM_BCM09_DP
  `undef DW_AXI_A2X_RM_BCM09_DP
`endif 

`ifdef DW_AXI_A2X_RM_BCM09_ECC
  `undef DW_AXI_A2X_RM_BCM09_ECC
`endif 

`ifdef DW_AXI_A2X_RM_BCM10
  `undef DW_AXI_A2X_RM_BCM10
`endif 

`ifdef DW_AXI_A2X_RM_BCM11
  `undef DW_AXI_A2X_RM_BCM11
`endif 

`ifdef DW_AXI_A2X_RM_BCM12
  `undef DW_AXI_A2X_RM_BCM12
`endif 

`ifdef DW_AXI_A2X_RM_BCM14
  `undef DW_AXI_A2X_RM_BCM14
`endif 

`ifdef DW_AXI_A2X_RM_BCM15
  `undef DW_AXI_A2X_RM_BCM15
`endif 

`ifdef DW_AXI_A2X_RM_BCM16
  `undef DW_AXI_A2X_RM_BCM16
`endif 

`ifdef DW_AXI_A2X_RM_BCM17
  `undef DW_AXI_A2X_RM_BCM17
`endif 

`ifdef DW_AXI_A2X_RM_BCM18_GEN
  `undef DW_AXI_A2X_RM_BCM18_GEN
`endif 

`ifdef DW_AXI_A2X_RM_BCM18_MON
  `undef DW_AXI_A2X_RM_BCM18_MON
`endif 

`ifdef DW_AXI_A2X_RM_BCM18_PGEN
  `undef DW_AXI_A2X_RM_BCM18_PGEN
`endif 

`ifdef DW_AXI_A2X_RM_BCM18_PGENA
  `undef DW_AXI_A2X_RM_BCM18_PGENA
`endif 

`ifdef DW_AXI_A2X_RM_BCM18_PMON
  `undef DW_AXI_A2X_RM_BCM18_PMON
`endif 

`ifdef DW_AXI_A2X_RM_BCM18_RS
  `undef DW_AXI_A2X_RM_BCM18_RS
`endif 

`ifdef DW_AXI_A2X_RM_BCM19_INTR
  `undef DW_AXI_A2X_RM_BCM19_INTR
`endif 

`ifdef DW_AXI_A2X_RM_BCM19_TRGT
  `undef DW_AXI_A2X_RM_BCM19_TRGT
`endif 

`ifdef DW_AXI_A2X_RM_BCM21
  `undef DW_AXI_A2X_RM_BCM21
`endif 

`ifdef DW_AXI_A2X_RM_BCM21_ATV
  `undef DW_AXI_A2X_RM_BCM21_ATV
`endif 

`ifdef DW_AXI_A2X_RM_BCM21_NEO
  `undef DW_AXI_A2X_RM_BCM21_NEO
`endif 

`ifdef DW_AXI_A2X_RM_BCM21_TGL
  `undef DW_AXI_A2X_RM_BCM21_TGL
`endif 

`ifdef DW_AXI_A2X_RM_BCM22
  `undef DW_AXI_A2X_RM_BCM22
`endif 

`ifdef DW_AXI_A2X_RM_BCM22_ATV
  `undef DW_AXI_A2X_RM_BCM22_ATV
`endif 

`ifdef DW_AXI_A2X_RM_BCM23
  `undef DW_AXI_A2X_RM_BCM23
`endif 

`ifdef DW_AXI_A2X_RM_BCM23_ATV
  `undef DW_AXI_A2X_RM_BCM23_ATV
`endif 

`ifdef DW_AXI_A2X_RM_BCM23_C
  `undef DW_AXI_A2X_RM_BCM23_C
`endif 

`ifdef DW_AXI_A2X_RM_BCM24
  `undef DW_AXI_A2X_RM_BCM24
`endif 

`ifdef DW_AXI_A2X_RM_BCM24_AP
  `undef DW_AXI_A2X_RM_BCM24_AP
`endif 

`ifdef DW_AXI_A2X_RM_BCM25
  `undef DW_AXI_A2X_RM_BCM25
`endif 

`ifdef DW_AXI_A2X_RM_BCM25_ATV
  `undef DW_AXI_A2X_RM_BCM25_ATV
`endif 

`ifdef DW_AXI_A2X_RM_BCM25_C
  `undef DW_AXI_A2X_RM_BCM25_C
`endif 

`ifdef DW_AXI_A2X_RM_BCM26
  `undef DW_AXI_A2X_RM_BCM26
`endif 

`ifdef DW_AXI_A2X_RM_BCM26_ATV
  `undef DW_AXI_A2X_RM_BCM26_ATV
`endif 

`ifdef DW_AXI_A2X_RM_BCM27
  `undef DW_AXI_A2X_RM_BCM27
`endif 

`ifdef DW_AXI_A2X_RM_BCM28
  `undef DW_AXI_A2X_RM_BCM28
`endif 

`ifdef DW_AXI_A2X_RM_BCM29
  `undef DW_AXI_A2X_RM_BCM29
`endif 

`ifdef DW_AXI_A2X_RM_BCM31_P2D_FIFOMEM
  `undef DW_AXI_A2X_RM_BCM31_P2D_FIFOMEM
`endif 

`ifdef DW_AXI_A2X_RM_BCM31_P2D_RD
  `undef DW_AXI_A2X_RM_BCM31_P2D_RD
`endif 

`ifdef DW_AXI_A2X_RM_BCM31_P2D_WR
  `undef DW_AXI_A2X_RM_BCM31_P2D_WR
`endif 

`ifdef DW_AXI_A2X_RM_BCM32_A
  `undef DW_AXI_A2X_RM_BCM32_A
`endif 

`ifdef DW_AXI_A2X_RM_BCM32_C
  `undef DW_AXI_A2X_RM_BCM32_C
`endif 

`ifdef DW_AXI_A2X_RM_BCM33_63_7_64_0
  `undef DW_AXI_A2X_RM_BCM33_63_7_64_0
`endif 

`ifdef DW_AXI_A2X_RM_BCM35
  `undef DW_AXI_A2X_RM_BCM35
`endif 

`ifdef DW_AXI_A2X_RM_BCM35_T
  `undef DW_AXI_A2X_RM_BCM35_T
`endif 

`ifdef DW_AXI_A2X_RM_BCM36
  `undef DW_AXI_A2X_RM_BCM36
`endif 

`ifdef DW_AXI_A2X_RM_BCM36_ACK
  `undef DW_AXI_A2X_RM_BCM36_ACK
`endif 

`ifdef DW_AXI_A2X_RM_BCM36_NHS
  `undef DW_AXI_A2X_RM_BCM36_NHS
`endif 

`ifdef DW_AXI_A2X_RM_BCM36_TGL
  `undef DW_AXI_A2X_RM_BCM36_TGL
`endif 

`ifdef DW_AXI_A2X_RM_BCM36_TGL_DO
  `undef DW_AXI_A2X_RM_BCM36_TGL_DO
`endif 

`ifdef DW_AXI_A2X_RM_BCM36_TGL_PLS
  `undef DW_AXI_A2X_RM_BCM36_TGL_PLS
`endif 

`ifdef DW_AXI_A2X_RM_BCM36_TGL_PLS_DO
  `undef DW_AXI_A2X_RM_BCM36_TGL_PLS_DO
`endif 

`ifdef DW_AXI_A2X_RM_BCM37
  `undef DW_AXI_A2X_RM_BCM37
`endif 

`ifdef DW_AXI_A2X_RM_BCM38
  `undef DW_AXI_A2X_RM_BCM38
`endif 

`ifdef DW_AXI_A2X_RM_BCM38_ADP
  `undef DW_AXI_A2X_RM_BCM38_ADP
`endif 

`ifdef DW_AXI_A2X_RM_BCM38_AP
  `undef DW_AXI_A2X_RM_BCM38_AP
`endif 

`ifdef DW_AXI_A2X_RM_BCM38_ECC
  `undef DW_AXI_A2X_RM_BCM38_ECC
`endif 

`ifdef DW_AXI_A2X_RM_BCM39
  `undef DW_AXI_A2X_RM_BCM39
`endif 

`ifdef DW_AXI_A2X_RM_BCM40
  `undef DW_AXI_A2X_RM_BCM40
`endif 

`ifdef DW_AXI_A2X_RM_BCM41
  `undef DW_AXI_A2X_RM_BCM41
`endif 

`ifdef DW_AXI_A2X_RM_BCM41_NEO
  `undef DW_AXI_A2X_RM_BCM41_NEO
`endif 

`ifdef DW_AXI_A2X_RM_BCM43
  `undef DW_AXI_A2X_RM_BCM43
`endif 

`ifdef DW_AXI_A2X_RM_BCM43_NRO
  `undef DW_AXI_A2X_RM_BCM43_NRO
`endif 

`ifdef DW_AXI_A2X_RM_BCM44
  `undef DW_AXI_A2X_RM_BCM44
`endif 

`ifdef DW_AXI_A2X_RM_BCM44_NRO
  `undef DW_AXI_A2X_RM_BCM44_NRO
`endif 

`ifdef DW_AXI_A2X_RM_BCM45_GN_D_A
  `undef DW_AXI_A2X_RM_BCM45_GN_D_A
`endif 

`ifdef DW_AXI_A2X_RM_BCM45_GN_D_AA
  `undef DW_AXI_A2X_RM_BCM45_GN_D_AA
`endif 

`ifdef DW_AXI_A2X_RM_BCM45_GN_D_B
  `undef DW_AXI_A2X_RM_BCM45_GN_D_B
`endif 

`ifdef DW_AXI_A2X_RM_BCM45_GN_D_C
  `undef DW_AXI_A2X_RM_BCM45_GN_D_C
`endif 

`ifdef DW_AXI_A2X_RM_BCM45_GN_D_D
  `undef DW_AXI_A2X_RM_BCM45_GN_D_D
`endif 

`ifdef DW_AXI_A2X_RM_BCM45_GN_D_E
  `undef DW_AXI_A2X_RM_BCM45_GN_D_E
`endif 

`ifdef DW_AXI_A2X_RM_BCM45_GN_D_F
  `undef DW_AXI_A2X_RM_BCM45_GN_D_F
`endif 

`ifdef DW_AXI_A2X_RM_BCM45_MN_D_A
  `undef DW_AXI_A2X_RM_BCM45_MN_D_A
`endif 

`ifdef DW_AXI_A2X_RM_BCM45_MN_D_AA
  `undef DW_AXI_A2X_RM_BCM45_MN_D_AA
`endif 

`ifdef DW_AXI_A2X_RM_BCM45_MN_D_B
  `undef DW_AXI_A2X_RM_BCM45_MN_D_B
`endif 

`ifdef DW_AXI_A2X_RM_BCM45_MN_D_C
  `undef DW_AXI_A2X_RM_BCM45_MN_D_C
`endif 

`ifdef DW_AXI_A2X_RM_BCM45_MN_D_D
  `undef DW_AXI_A2X_RM_BCM45_MN_D_D
`endif 

`ifdef DW_AXI_A2X_RM_BCM45_MN_D_E
  `undef DW_AXI_A2X_RM_BCM45_MN_D_E
`endif 

`ifdef DW_AXI_A2X_RM_BCM45_MN_D_F
  `undef DW_AXI_A2X_RM_BCM45_MN_D_F
`endif 

`ifdef DW_AXI_A2X_RM_BCM46_A
  `undef DW_AXI_A2X_RM_BCM46_A
`endif 

`ifdef DW_AXI_A2X_RM_BCM46_AA
  `undef DW_AXI_A2X_RM_BCM46_AA
`endif 

`ifdef DW_AXI_A2X_RM_BCM46_B
  `undef DW_AXI_A2X_RM_BCM46_B
`endif 

`ifdef DW_AXI_A2X_RM_BCM46_B_32A
  `undef DW_AXI_A2X_RM_BCM46_B_32A
`endif 

`ifdef DW_AXI_A2X_RM_BCM46_C
  `undef DW_AXI_A2X_RM_BCM46_C
`endif 

`ifdef DW_AXI_A2X_RM_BCM46_C_64A
  `undef DW_AXI_A2X_RM_BCM46_C_64A
`endif 

`ifdef DW_AXI_A2X_RM_BCM46_D
  `undef DW_AXI_A2X_RM_BCM46_D
`endif 

`ifdef DW_AXI_A2X_RM_BCM46_D_128A
  `undef DW_AXI_A2X_RM_BCM46_D_128A
`endif 

`ifdef DW_AXI_A2X_RM_BCM46_E
  `undef DW_AXI_A2X_RM_BCM46_E
`endif 

`ifdef DW_AXI_A2X_RM_BCM46_F
  `undef DW_AXI_A2X_RM_BCM46_F
`endif 

`ifdef DW_AXI_A2X_RM_BCM46_X
  `undef DW_AXI_A2X_RM_BCM46_X
`endif 

`ifdef DW_AXI_A2X_RM_BCM47
  `undef DW_AXI_A2X_RM_BCM47
`endif 

`ifdef DW_AXI_A2X_RM_BCM48
  `undef DW_AXI_A2X_RM_BCM48
`endif 

`ifdef DW_AXI_A2X_RM_BCM48_DM
  `undef DW_AXI_A2X_RM_BCM48_DM
`endif 

`ifdef DW_AXI_A2X_RM_BCM48_SV
  `undef DW_AXI_A2X_RM_BCM48_SV
`endif 

`ifdef DW_AXI_A2X_RM_BCM49
  `undef DW_AXI_A2X_RM_BCM49
`endif 

`ifdef DW_AXI_A2X_RM_BCM49_SV
  `undef DW_AXI_A2X_RM_BCM49_SV
`endif 

`ifdef DW_AXI_A2X_RM_BCM50
  `undef DW_AXI_A2X_RM_BCM50
`endif 

`ifdef DW_AXI_A2X_RM_BCM51
  `undef DW_AXI_A2X_RM_BCM51
`endif 

`ifdef DW_AXI_A2X_RM_BCM52
  `undef DW_AXI_A2X_RM_BCM52
`endif 

`ifdef DW_AXI_A2X_RM_BCM53
  `undef DW_AXI_A2X_RM_BCM53
`endif 

`ifdef DW_AXI_A2X_RM_BCM54
  `undef DW_AXI_A2X_RM_BCM54
`endif 

`ifdef DW_AXI_A2X_RM_BCM55
  `undef DW_AXI_A2X_RM_BCM55
`endif 

`ifdef DW_AXI_A2X_RM_BCM55_C
  `undef DW_AXI_A2X_RM_BCM55_C
`endif 

`ifdef DW_AXI_A2X_RM_BCM56
  `undef DW_AXI_A2X_RM_BCM56
`endif 

`ifdef DW_AXI_A2X_RM_BCM57
  `undef DW_AXI_A2X_RM_BCM57
`endif 

`ifdef DW_AXI_A2X_RM_BCM57_ATV
  `undef DW_AXI_A2X_RM_BCM57_ATV
`endif 

`ifdef DW_AXI_A2X_RM_BCM58
  `undef DW_AXI_A2X_RM_BCM58
`endif 

`ifdef DW_AXI_A2X_RM_BCM58_ATV
  `undef DW_AXI_A2X_RM_BCM58_ATV
`endif 

`ifdef DW_AXI_A2X_RM_BCM59
  `undef DW_AXI_A2X_RM_BCM59
`endif 

`ifdef DW_AXI_A2X_RM_BCM60
  `undef DW_AXI_A2X_RM_BCM60
`endif 

`ifdef DW_AXI_A2X_RM_BCM62
  `undef DW_AXI_A2X_RM_BCM62
`endif 

`ifdef DW_AXI_A2X_RM_BCM63
  `undef DW_AXI_A2X_RM_BCM63
`endif 

`ifdef DW_AXI_A2X_RM_BCM64
  `undef DW_AXI_A2X_RM_BCM64
`endif 

`ifdef DW_AXI_A2X_RM_BCM64_TD
  `undef DW_AXI_A2X_RM_BCM64_TD
`endif 

`ifdef DW_AXI_A2X_RM_BCM65
  `undef DW_AXI_A2X_RM_BCM65
`endif 

`ifdef DW_AXI_A2X_RM_BCM65_ATV
  `undef DW_AXI_A2X_RM_BCM65_ATV
`endif 

`ifdef DW_AXI_A2X_RM_BCM65_TD
  `undef DW_AXI_A2X_RM_BCM65_TD
`endif 

`ifdef DW_AXI_A2X_RM_BCM66
  `undef DW_AXI_A2X_RM_BCM66
`endif 

`ifdef DW_AXI_A2X_RM_BCM66_ATV
  `undef DW_AXI_A2X_RM_BCM66_ATV
`endif 

`ifdef DW_AXI_A2X_RM_BCM66_DMS
  `undef DW_AXI_A2X_RM_BCM66_DMS
`endif 

`ifdef DW_AXI_A2X_RM_BCM66_DMS_ATV
  `undef DW_AXI_A2X_RM_BCM66_DMS_ATV
`endif 

`ifdef DW_AXI_A2X_RM_BCM66_EFES
  `undef DW_AXI_A2X_RM_BCM66_EFES
`endif 

`ifdef DW_AXI_A2X_RM_BCM66_PR
  `undef DW_AXI_A2X_RM_BCM66_PR
`endif 

`ifdef DW_AXI_A2X_RM_BCM66_WAE
  `undef DW_AXI_A2X_RM_BCM66_WAE
`endif 

`ifdef DW_AXI_A2X_RM_BCM66_WAE_ATV
  `undef DW_AXI_A2X_RM_BCM66_WAE_ATV
`endif 

`ifdef DW_AXI_A2X_RM_BCM68_63_7_0
  `undef DW_AXI_A2X_RM_BCM68_63_7_0
`endif 

`ifdef DW_AXI_A2X_RM_BCM69_63_7_0
  `undef DW_AXI_A2X_RM_BCM69_63_7_0
`endif 

`ifdef DW_AXI_A2X_RM_BCM70_63_7_0_0
  `undef DW_AXI_A2X_RM_BCM70_63_7_0_0
`endif 

`ifdef DW_AXI_A2X_RM_BCM71
  `undef DW_AXI_A2X_RM_BCM71
`endif 

`ifdef DW_AXI_A2X_RM_BCM72
  `undef DW_AXI_A2X_RM_BCM72
`endif 

`ifdef DW_AXI_A2X_RM_BCM74
  `undef DW_AXI_A2X_RM_BCM74
`endif 

`ifdef DW_AXI_A2X_RM_BCM76
  `undef DW_AXI_A2X_RM_BCM76
`endif 

`ifdef DW_AXI_A2X_RM_BCM77
  `undef DW_AXI_A2X_RM_BCM77
`endif 

`ifdef DW_AXI_A2X_RM_BCM78
  `undef DW_AXI_A2X_RM_BCM78
`endif 

`ifdef DW_AXI_A2X_RM_BCM79
  `undef DW_AXI_A2X_RM_BCM79
`endif 

`ifdef DW_AXI_A2X_RM_BCM79_MO
  `undef DW_AXI_A2X_RM_BCM79_MO
`endif 

`ifdef DW_AXI_A2X_RM_BCM83_GEN
  `undef DW_AXI_A2X_RM_BCM83_GEN
`endif 

`ifdef DW_AXI_A2X_RM_BCM84_MON
  `undef DW_AXI_A2X_RM_BCM84_MON
`endif 

`ifdef DW_AXI_A2X_RM_BCM85
  `undef DW_AXI_A2X_RM_BCM85
`endif 

`ifdef DW_AXI_A2X_RM_BCM86
  `undef DW_AXI_A2X_RM_BCM86
`endif 

`ifdef DW_AXI_A2X_RM_BCM87
  `undef DW_AXI_A2X_RM_BCM87
`endif 

`ifdef DW_AXI_A2X_RM_BCM90
  `undef DW_AXI_A2X_RM_BCM90
`endif 

`ifdef DW_AXI_A2X_RM_BCM91
  `undef DW_AXI_A2X_RM_BCM91
`endif 

`ifdef DW_AXI_A2X_RM_BCM92
  `undef DW_AXI_A2X_RM_BCM92
`endif 

`ifdef DW_AXI_A2X_RM_BCM92_AD
  `undef DW_AXI_A2X_RM_BCM92_AD
`endif 

`ifdef DW_AXI_A2X_RM_BCM92_AD_DO
  `undef DW_AXI_A2X_RM_BCM92_AD_DO
`endif 

`ifdef DW_AXI_A2X_RM_BCM92_RD
  `undef DW_AXI_A2X_RM_BCM92_RD
`endif 

`ifdef DW_AXI_A2X_RM_BCM92_RD_AD
  `undef DW_AXI_A2X_RM_BCM92_RD_AD
`endif 

`ifdef DW_AXI_A2X_RM_BCM92_RD_AD_DO
  `undef DW_AXI_A2X_RM_BCM92_RD_AD_DO
`endif 

`ifdef DW_AXI_A2X_RM_BCM92_RD_DO
  `undef DW_AXI_A2X_RM_BCM92_RD_DO
`endif 

`ifdef DW_AXI_A2X_RM_BCM93
  `undef DW_AXI_A2X_RM_BCM93
`endif 

`ifdef DW_AXI_A2X_RM_BCM93_NDSVA
  `undef DW_AXI_A2X_RM_BCM93_NDSVA
`endif 

`ifdef DW_AXI_A2X_RM_BCM94
  `undef DW_AXI_A2X_RM_BCM94
`endif 

`ifdef DW_AXI_A2X_RM_BCM95
  `undef DW_AXI_A2X_RM_BCM95
`endif 

`ifdef DW_AXI_A2X_RM_BCM95_E
  `undef DW_AXI_A2X_RM_BCM95_E
`endif 

`ifdef DW_AXI_A2X_RM_BCM95_I
  `undef DW_AXI_A2X_RM_BCM95_I
`endif 

`ifdef DW_AXI_A2X_RM_BCM95_IE
  `undef DW_AXI_A2X_RM_BCM95_IE
`endif 

`ifdef DW_AXI_A2X_RM_BCM95_NE
  `undef DW_AXI_A2X_RM_BCM95_NE
`endif 

`ifdef DW_AXI_A2X_RM_BCM95_NE_E
  `undef DW_AXI_A2X_RM_BCM95_NE_E
`endif 

`ifdef DW_AXI_A2X_RM_BCM95_NE_I
  `undef DW_AXI_A2X_RM_BCM95_NE_I
`endif 

`ifdef DW_AXI_A2X_RM_BCM95_NE_IE
  `undef DW_AXI_A2X_RM_BCM95_NE_IE
`endif 

`ifdef DW_AXI_A2X_RM_BCM98
  `undef DW_AXI_A2X_RM_BCM98
`endif 

`ifdef DW_AXI_A2X_RM_BCM99
  `undef DW_AXI_A2X_RM_BCM99
`endif 

`ifdef DW_AXI_A2X_RM_BCM99_3
  `undef DW_AXI_A2X_RM_BCM99_3
`endif 

`ifdef DW_AXI_A2X_RM_BCM99_4
  `undef DW_AXI_A2X_RM_BCM99_4
`endif 

`ifdef DW_AXI_A2X_RM_BCM99_N
  `undef DW_AXI_A2X_RM_BCM99_N
`endif 

`ifdef DW_AXI_A2X_RM_BVM01
  `undef DW_AXI_A2X_RM_BVM01
`endif 

`ifdef DW_AXI_A2X_RM_BVM02
  `undef DW_AXI_A2X_RM_BVM02
`endif 

`ifdef DW_AXI_A2X_RM_SVA01
  `undef DW_AXI_A2X_RM_SVA01
`endif 

`ifdef DW_AXI_A2X_RM_SVA02
  `undef DW_AXI_A2X_RM_SVA02
`endif 

`ifdef DW_AXI_A2X_RM_SVA03
  `undef DW_AXI_A2X_RM_SVA03
`endif 

`ifdef DW_AXI_A2X_RM_SVA04
  `undef DW_AXI_A2X_RM_SVA04
`endif 

`ifdef DW_AXI_A2X_RM_SVA05
  `undef DW_AXI_A2X_RM_SVA05
`endif 

`ifdef DW_AXI_A2X_RM_SVA06
  `undef DW_AXI_A2X_RM_SVA06
`endif 

`ifdef DW_AXI_A2X_RM_SVA07
  `undef DW_AXI_A2X_RM_SVA07
`endif 

`ifdef DW_AXI_A2X_RM_SVA08
  `undef DW_AXI_A2X_RM_SVA08
`endif 

`ifdef DW_AXI_A2X_RM_SVA09
  `undef DW_AXI_A2X_RM_SVA09
`endif 

`ifdef DW_AXI_A2X_RM_SVA10
  `undef DW_AXI_A2X_RM_SVA10
`endif 

`ifdef DW_AXI_A2X_RM_SVA11
  `undef DW_AXI_A2X_RM_SVA11
`endif 

`ifdef DW_AXI_A2X_RM_SVA12_A
  `undef DW_AXI_A2X_RM_SVA12_A
`endif 

`ifdef DW_AXI_A2X_RM_SVA12_B
  `undef DW_AXI_A2X_RM_SVA12_B
`endif 

`ifdef DW_AXI_A2X_RM_SVA12_C
  `undef DW_AXI_A2X_RM_SVA12_C
`endif 

`ifdef DW_AXI_A2X_RM_SVA99
  `undef DW_AXI_A2X_RM_SVA99
`endif 

`ifdef __GUARD__DW_AXI_A2X_ALL_INCLUDES__VH__
  `undef __GUARD__DW_AXI_A2X_ALL_INCLUDES__VH__
`endif 

`ifdef cb_dummy_parameter_definition
  `undef cb_dummy_parameter_definition
`endif 

