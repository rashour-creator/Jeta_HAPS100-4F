//##########################################################
// Generated unprefix file for workspace: DW_axi_a2x
//##########################################################

`ifdef i_axi_a2x_2___GUARD__DW_AXI_A2X_DEFINE_CONSTANTS__VH__
  `define __GUARD__DW_AXI_A2X_DEFINE_CONSTANTS__VH__ `i_axi_a2x_2___GUARD__DW_AXI_A2X_DEFINE_CONSTANTS__VH__
`endif 

`ifdef i_axi_a2x_2_A2X_BSW
  `define A2X_BSW `i_axi_a2x_2_A2X_BSW
`endif 

`ifdef i_axi_a2x_2_A2X_BTW
  `define A2X_BTW `i_axi_a2x_2_A2X_BTW
`endif 

`ifdef i_axi_a2x_2_A2X_LTW
  `define A2X_LTW `i_axi_a2x_2_A2X_LTW
`endif 

`ifdef i_axi_a2x_2_A2X_CTW
  `define A2X_CTW `i_axi_a2x_2_A2X_CTW
`endif 

`ifdef i_axi_a2x_2_A2X_PTW
  `define A2X_PTW `i_axi_a2x_2_A2X_PTW
`endif 

`ifdef i_axi_a2x_2_A2X_RSW
  `define A2X_RSW `i_axi_a2x_2_A2X_RSW
`endif 

`ifdef i_axi_a2x_2_A2X_BRESPW
  `define A2X_BRESPW `i_axi_a2x_2_A2X_BRESPW
`endif 

`ifdef i_axi_a2x_2_A2X_RRESPW
  `define A2X_RRESPW `i_axi_a2x_2_A2X_RRESPW
`endif 

`ifdef i_axi_a2x_2_A2X_HIDW
  `define A2X_HIDW `i_axi_a2x_2_A2X_HIDW
`endif 

`ifdef i_axi_a2x_2_A2X_HBLW
  `define A2X_HBLW `i_axi_a2x_2_A2X_HBLW
`endif 

`ifdef i_axi_a2x_2_A2X_HBTYPE_W
  `define A2X_HBTYPE_W `i_axi_a2x_2_A2X_HBTYPE_W
`endif 

`ifdef i_axi_a2x_2_A2X_MAX_BSBW
  `define A2X_MAX_BSBW `i_axi_a2x_2_A2X_MAX_BSBW
`endif 

`ifdef i_axi_a2x_2_CT_MODE
  `define CT_MODE `i_axi_a2x_2_CT_MODE
`endif 

`ifdef i_axi_a2x_2_SNF_MODE
  `define SNF_MODE `i_axi_a2x_2_SNF_MODE
`endif 

`ifdef i_axi_a2x_2_ABURST_FIXED
  `define ABURST_FIXED `i_axi_a2x_2_ABURST_FIXED
`endif 

`ifdef i_axi_a2x_2_ABURST_INCR
  `define ABURST_INCR `i_axi_a2x_2_ABURST_INCR
`endif 

`ifdef i_axi_a2x_2_ABURST_WRAP
  `define ABURST_WRAP `i_axi_a2x_2_ABURST_WRAP
`endif 

`ifdef i_axi_a2x_2_HTRANS_IDLE
  `define HTRANS_IDLE `i_axi_a2x_2_HTRANS_IDLE
`endif 

`ifdef i_axi_a2x_2_HTRANS_BUSY
  `define HTRANS_BUSY `i_axi_a2x_2_HTRANS_BUSY
`endif 

`ifdef i_axi_a2x_2_HTRANS_NSEQ
  `define HTRANS_NSEQ `i_axi_a2x_2_HTRANS_NSEQ
`endif 

`ifdef i_axi_a2x_2_HTRANS_SEQ
  `define HTRANS_SEQ `i_axi_a2x_2_HTRANS_SEQ
`endif 

`ifdef i_axi_a2x_2_HBURST_SINGLE
  `define HBURST_SINGLE `i_axi_a2x_2_HBURST_SINGLE
`endif 

`ifdef i_axi_a2x_2_HBURST_INCR
  `define HBURST_INCR `i_axi_a2x_2_HBURST_INCR
`endif 

`ifdef i_axi_a2x_2_HBURST_WRAP4
  `define HBURST_WRAP4 `i_axi_a2x_2_HBURST_WRAP4
`endif 

`ifdef i_axi_a2x_2_HBURST_INCR4
  `define HBURST_INCR4 `i_axi_a2x_2_HBURST_INCR4
`endif 

`ifdef i_axi_a2x_2_HBURST_WRAP8
  `define HBURST_WRAP8 `i_axi_a2x_2_HBURST_WRAP8
`endif 

`ifdef i_axi_a2x_2_HBURST_INCR8
  `define HBURST_INCR8 `i_axi_a2x_2_HBURST_INCR8
`endif 

`ifdef i_axi_a2x_2_HBURST_WRAP16
  `define HBURST_WRAP16 `i_axi_a2x_2_HBURST_WRAP16
`endif 

`ifdef i_axi_a2x_2_HBURST_INCR16
  `define HBURST_INCR16 `i_axi_a2x_2_HBURST_INCR16
`endif 

`ifdef i_axi_a2x_2_HSIZE_8
  `define HSIZE_8 `i_axi_a2x_2_HSIZE_8
`endif 

`ifdef i_axi_a2x_2_HSIZE_16
  `define HSIZE_16 `i_axi_a2x_2_HSIZE_16
`endif 

`ifdef i_axi_a2x_2_HSIZE_32
  `define HSIZE_32 `i_axi_a2x_2_HSIZE_32
`endif 

`ifdef i_axi_a2x_2_HSIZE_64
  `define HSIZE_64 `i_axi_a2x_2_HSIZE_64
`endif 

`ifdef i_axi_a2x_2_HSIZE_128
  `define HSIZE_128 `i_axi_a2x_2_HSIZE_128
`endif 

`ifdef i_axi_a2x_2_HSIZE_256
  `define HSIZE_256 `i_axi_a2x_2_HSIZE_256
`endif 

`ifdef i_axi_a2x_2_HSIZE_512
  `define HSIZE_512 `i_axi_a2x_2_HSIZE_512
`endif 

`ifdef i_axi_a2x_2_HSIZE_1024
  `define HSIZE_1024 `i_axi_a2x_2_HSIZE_1024
`endif 

`ifdef i_axi_a2x_2_HSIZE_8BIT
  `define HSIZE_8BIT `i_axi_a2x_2_HSIZE_8BIT
`endif 

`ifdef i_axi_a2x_2_HSIZE_16BIT
  `define HSIZE_16BIT `i_axi_a2x_2_HSIZE_16BIT
`endif 

`ifdef i_axi_a2x_2_HSIZE_32BIT
  `define HSIZE_32BIT `i_axi_a2x_2_HSIZE_32BIT
`endif 

`ifdef i_axi_a2x_2_HSIZE_64BIT
  `define HSIZE_64BIT `i_axi_a2x_2_HSIZE_64BIT
`endif 

`ifdef i_axi_a2x_2_HSIZE_128BIT
  `define HSIZE_128BIT `i_axi_a2x_2_HSIZE_128BIT
`endif 

`ifdef i_axi_a2x_2_HSIZE_256BIT
  `define HSIZE_256BIT `i_axi_a2x_2_HSIZE_256BIT
`endif 

`ifdef i_axi_a2x_2_HSIZE_512BIT
  `define HSIZE_512BIT `i_axi_a2x_2_HSIZE_512BIT
`endif 

`ifdef i_axi_a2x_2_HSIZE_1024BIT
  `define HSIZE_1024BIT `i_axi_a2x_2_HSIZE_1024BIT
`endif 

`ifdef i_axi_a2x_2_HSIZE_BYTE
  `define HSIZE_BYTE `i_axi_a2x_2_HSIZE_BYTE
`endif 

`ifdef i_axi_a2x_2_HSIZE_WORD16
  `define HSIZE_WORD16 `i_axi_a2x_2_HSIZE_WORD16
`endif 

`ifdef i_axi_a2x_2_HSIZE_WORD32
  `define HSIZE_WORD32 `i_axi_a2x_2_HSIZE_WORD32
`endif 

`ifdef i_axi_a2x_2_HSIZE_WORD64
  `define HSIZE_WORD64 `i_axi_a2x_2_HSIZE_WORD64
`endif 

`ifdef i_axi_a2x_2_HSIZE_WORD128
  `define HSIZE_WORD128 `i_axi_a2x_2_HSIZE_WORD128
`endif 

`ifdef i_axi_a2x_2_HSIZE_WORD256
  `define HSIZE_WORD256 `i_axi_a2x_2_HSIZE_WORD256
`endif 

`ifdef i_axi_a2x_2_HSIZE_WORD512
  `define HSIZE_WORD512 `i_axi_a2x_2_HSIZE_WORD512
`endif 

`ifdef i_axi_a2x_2_HSIZE_WORD1024
  `define HSIZE_WORD1024 `i_axi_a2x_2_HSIZE_WORD1024
`endif 

`ifdef i_axi_a2x_2_HPROT_DATA
  `define HPROT_DATA `i_axi_a2x_2_HPROT_DATA
`endif 

`ifdef i_axi_a2x_2_HPROT_PRIV
  `define HPROT_PRIV `i_axi_a2x_2_HPROT_PRIV
`endif 

`ifdef i_axi_a2x_2_HPROT_BUFF
  `define HPROT_BUFF `i_axi_a2x_2_HPROT_BUFF
`endif 

`ifdef i_axi_a2x_2_HPROT_CACHE
  `define HPROT_CACHE `i_axi_a2x_2_HPROT_CACHE
`endif 

`ifdef i_axi_a2x_2_HRESP_OKAY
  `define HRESP_OKAY `i_axi_a2x_2_HRESP_OKAY
`endif 

`ifdef i_axi_a2x_2_HRESP_ERROR
  `define HRESP_ERROR `i_axi_a2x_2_HRESP_ERROR
`endif 

`ifdef i_axi_a2x_2_HRESP_RETRY
  `define HRESP_RETRY `i_axi_a2x_2_HRESP_RETRY
`endif 

`ifdef i_axi_a2x_2_HRESP_SPLIT
  `define HRESP_SPLIT `i_axi_a2x_2_HRESP_SPLIT
`endif 

`ifdef i_axi_a2x_2_AFIXED
  `define AFIXED `i_axi_a2x_2_AFIXED
`endif 

`ifdef i_axi_a2x_2_AINCR
  `define AINCR `i_axi_a2x_2_AINCR
`endif 

`ifdef i_axi_a2x_2_AWRAP
  `define AWRAP `i_axi_a2x_2_AWRAP
`endif 

`ifdef i_axi_a2x_2_AOKAY
  `define AOKAY `i_axi_a2x_2_AOKAY
`endif 

`ifdef i_axi_a2x_2_AEXOKAY
  `define AEXOKAY `i_axi_a2x_2_AEXOKAY
`endif 

`ifdef i_axi_a2x_2_ASLVERR
  `define ASLVERR `i_axi_a2x_2_ASLVERR
`endif 

`ifdef i_axi_a2x_2_ADECERR
  `define ADECERR `i_axi_a2x_2_ADECERR
`endif 

`ifdef i_axi_a2x_2___GUARD__DW_AXI_A2X_CC_CONSTANTS__VH__
  `define __GUARD__DW_AXI_A2X_CC_CONSTANTS__VH__ `i_axi_a2x_2___GUARD__DW_AXI_A2X_CC_CONSTANTS__VH__
`endif 

`ifdef i_axi_a2x_2_USE_FOUNDATION
  `define USE_FOUNDATION `i_axi_a2x_2_USE_FOUNDATION
`endif 

`ifdef i_axi_a2x_2_A2X_USE_FOUNDATION
  `define A2X_USE_FOUNDATION `i_axi_a2x_2_A2X_USE_FOUNDATION
`endif 

`ifdef i_axi_a2x_2_A2X_LOWPWR_IF
  `define A2X_LOWPWR_IF `i_axi_a2x_2_A2X_LOWPWR_IF
`endif 

`ifdef i_axi_a2x_2_A2X_LOWPWR_NOPX_CNT
  `define A2X_LOWPWR_NOPX_CNT `i_axi_a2x_2_A2X_LOWPWR_NOPX_CNT
`endif 

`ifdef i_axi_a2x_2_A2X_PP_MODE
  `define A2X_PP_MODE `i_axi_a2x_2_A2X_PP_MODE
`endif 

`ifdef i_axi_a2x_2_A2X_AHB_INTERFACE_TYPE
  `define A2X_AHB_INTERFACE_TYPE `i_axi_a2x_2_A2X_AHB_INTERFACE_TYPE
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_EXTD_MEMTYPE
  `define A2X_HAS_EXTD_MEMTYPE `i_axi_a2x_2_A2X_HAS_EXTD_MEMTYPE
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_SECURE_XFER
  `define A2X_HAS_SECURE_XFER `i_axi_a2x_2_A2X_HAS_SECURE_XFER
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_EXCL_XFER
  `define A2X_HAS_EXCL_XFER `i_axi_a2x_2_A2X_HAS_EXCL_XFER
`endif 

`ifdef i_axi_a2x_2_A2X_HPTW
  `define A2X_HPTW `i_axi_a2x_2_A2X_HPTW
`endif 

`ifdef i_axi_a2x_2_A2X_AXI_INTERFACE_TYPE
  `define A2X_AXI_INTERFACE_TYPE `i_axi_a2x_2_A2X_AXI_INTERFACE_TYPE
`endif 

`ifdef i_axi_a2x_2_A2X_INT_AXI3
  `define A2X_INT_AXI3 `i_axi_a2x_2_A2X_INT_AXI3
`endif 

`ifdef i_axi_a2x_2_A2X_INT_LTW
  `define A2X_INT_LTW `i_axi_a2x_2_A2X_INT_LTW
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_AXI3
  `define A2X_HAS_AXI3 `i_axi_a2x_2_A2X_HAS_AXI3
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_AXI4
  `define A2X_HAS_AXI4 `i_axi_a2x_2_A2X_HAS_AXI4
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_ACELITE
  `define A2X_HAS_ACELITE `i_axi_a2x_2_A2X_HAS_ACELITE
`endif 

`ifdef i_axi_a2x_2_A2X_AHB_LITE_MODE
  `define A2X_AHB_LITE_MODE `i_axi_a2x_2_A2X_AHB_LITE_MODE
`endif 

`ifdef i_axi_a2x_2_A2X_AHB_SCALAR_HRESP
  `define A2X_AHB_SCALAR_HRESP `i_axi_a2x_2_A2X_AHB_SCALAR_HRESP
`endif 

`ifdef i_axi_a2x_2_A2X_AHB_SPLIT_MODE
  `define A2X_AHB_SPLIT_MODE `i_axi_a2x_2_A2X_AHB_SPLIT_MODE
`endif 

`ifdef i_axi_a2x_2_AHB_SPLIT_MODE
  `define AHB_SPLIT_MODE `i_axi_a2x_2_AHB_SPLIT_MODE
`endif 

`ifdef i_axi_a2x_2_A2X_NUM_AHBM
  `define A2X_NUM_AHBM `i_axi_a2x_2_A2X_NUM_AHBM
`endif 

`ifdef i_axi_a2x_2_A2X_HREADY_LOW_PERIOD
  `define A2X_HREADY_LOW_PERIOD `i_axi_a2x_2_A2X_HREADY_LOW_PERIOD
`endif 

`ifdef i_axi_a2x_2_A2X_LOCKED
  `define A2X_LOCKED `i_axi_a2x_2_A2X_LOCKED
`endif 

`ifdef i_axi_a2x_2_A2X_CLK_MODE
  `define A2X_CLK_MODE `i_axi_a2x_2_A2X_CLK_MODE
`endif 

`ifdef i_axi_a2x_2_A2X_PP_SYNC_DEPTH
  `define A2X_PP_SYNC_DEPTH `i_axi_a2x_2_A2X_PP_SYNC_DEPTH
`endif 

`ifdef i_axi_a2x_2_F_SYNC_TYPE_PP
  `define F_SYNC_TYPE_PP `i_axi_a2x_2_F_SYNC_TYPE_PP
`endif 

`ifdef i_axi_a2x_2_A2X_SP_SYNC_DEPTH
  `define A2X_SP_SYNC_DEPTH `i_axi_a2x_2_A2X_SP_SYNC_DEPTH
`endif 

`ifdef i_axi_a2x_2_F_SYNC_TYPE_SP
  `define F_SYNC_TYPE_SP `i_axi_a2x_2_F_SYNC_TYPE_SP
`endif 

`ifdef i_axi_a2x_2_A2X_SYNC_DEPTH_BUSY
  `define A2X_SYNC_DEPTH_BUSY `i_axi_a2x_2_A2X_SYNC_DEPTH_BUSY
`endif 

`ifdef i_axi_a2x_2_A2X_PP_IDW
  `define A2X_PP_IDW `i_axi_a2x_2_A2X_PP_IDW
`endif 

`ifdef i_axi_a2x_2_A2X_IDW
  `define A2X_IDW `i_axi_a2x_2_A2X_IDW
`endif 

`ifdef i_axi_a2x_2_A2X_SP_IDW
  `define A2X_SP_IDW `i_axi_a2x_2_A2X_SP_IDW
`endif 

`ifdef i_axi_a2x_2_A2X_PP_AW
  `define A2X_PP_AW `i_axi_a2x_2_A2X_PP_AW
`endif 

`ifdef i_axi_a2x_2_A2X_AW
  `define A2X_AW `i_axi_a2x_2_A2X_AW
`endif 

`ifdef i_axi_a2x_2_A2X_SP_AW
  `define A2X_SP_AW `i_axi_a2x_2_A2X_SP_AW
`endif 

`ifdef i_axi_a2x_2_A2X_BOUNDARY_W
  `define A2X_BOUNDARY_W `i_axi_a2x_2_A2X_BOUNDARY_W
`endif 

`ifdef i_axi_a2x_2_A2X_PP_BLW
  `define A2X_PP_BLW `i_axi_a2x_2_A2X_PP_BLW
`endif 

`ifdef i_axi_a2x_2_A2X_SP_BLW
  `define A2X_SP_BLW `i_axi_a2x_2_A2X_SP_BLW
`endif 

`ifdef i_axi_a2x_2_A2X_BLW
  `define A2X_BLW `i_axi_a2x_2_A2X_BLW
`endif 

`ifdef i_axi_a2x_2_A2X_MAX_ALEN
  `define A2X_MAX_ALEN `i_axi_a2x_2_A2X_MAX_ALEN
`endif 

`ifdef i_axi_a2x_2_A2X_PP_DW
  `define A2X_PP_DW `i_axi_a2x_2_A2X_PP_DW
`endif 

`ifdef i_axi_a2x_2_A2X_SP_DW
  `define A2X_SP_DW `i_axi_a2x_2_A2X_SP_DW
`endif 

`ifdef i_axi_a2x_2_A2X_RS_RATIO
  `define A2X_RS_RATIO `i_axi_a2x_2_A2X_RS_RATIO
`endif 

`ifdef i_axi_a2x_2_A2X_RS_RATIO_LOG2
  `define A2X_RS_RATIO_LOG2 `i_axi_a2x_2_A2X_RS_RATIO_LOG2
`endif 

`ifdef i_axi_a2x_2_A2X_PP_ENDIAN
  `define A2X_PP_ENDIAN `i_axi_a2x_2_A2X_PP_ENDIAN
`endif 

`ifdef i_axi_a2x_2_A2X_SP_ENDIAN
  `define A2X_SP_ENDIAN `i_axi_a2x_2_A2X_SP_ENDIAN
`endif 

`ifdef i_axi_a2x_2_A2X_WBUF_MODE
  `define A2X_WBUF_MODE `i_axi_a2x_2_A2X_WBUF_MODE
`endif 

`ifdef i_axi_a2x_2_A2X_HCBUF_MODE
  `define A2X_HCBUF_MODE `i_axi_a2x_2_A2X_HCBUF_MODE
`endif 

`ifdef i_axi_a2x_2_A2X_APB_MODE
  `define A2X_APB_MODE `i_axi_a2x_2_A2X_APB_MODE
`endif 

`ifdef i_axi_a2x_2_A2X_HCSNF_WLEN
  `define A2X_HCSNF_WLEN `i_axi_a2x_2_A2X_HCSNF_WLEN
`endif 

`ifdef i_axi_a2x_2_A2X_SNF_AWLEN_DFLT
  `define A2X_SNF_AWLEN_DFLT `i_axi_a2x_2_A2X_SNF_AWLEN_DFLT
`endif 

`ifdef i_axi_a2x_2_A2X_SNF_AWLEN_MIN
  `define A2X_SNF_AWLEN_MIN `i_axi_a2x_2_A2X_SNF_AWLEN_MIN
`endif 

`ifdef i_axi_a2x_2_A2X_HINCR_HCBCNT
  `define A2X_HINCR_HCBCNT `i_axi_a2x_2_A2X_HINCR_HCBCNT
`endif 

`ifdef i_axi_a2x_2_A2X_SINGLE_RBCNT
  `define A2X_SINGLE_RBCNT `i_axi_a2x_2_A2X_SINGLE_RBCNT
`endif 

`ifdef i_axi_a2x_2_A2X_SINGLE_WBCNT
  `define A2X_SINGLE_WBCNT `i_axi_a2x_2_A2X_SINGLE_WBCNT
`endif 

`ifdef i_axi_a2x_2_A2X_HINCR_WBCNT_MIN
  `define A2X_HINCR_WBCNT_MIN `i_axi_a2x_2_A2X_HINCR_WBCNT_MIN
`endif 

`ifdef i_axi_a2x_2_A2X_HINCR_WBCNT_MAX
  `define A2X_HINCR_WBCNT_MAX `i_axi_a2x_2_A2X_HINCR_WBCNT_MAX
`endif 

`ifdef i_axi_a2x_2_A2X_HINCR_AWLEN_DFLT
  `define A2X_HINCR_AWLEN_DFLT `i_axi_a2x_2_A2X_HINCR_AWLEN_DFLT
`endif 

`ifdef i_axi_a2x_2_A2X_HINCR_AWLEN_MIN
  `define A2X_HINCR_AWLEN_MIN `i_axi_a2x_2_A2X_HINCR_AWLEN_MIN
`endif 

`ifdef i_axi_a2x_2_A2X_BRESP_MODE
  `define A2X_BRESP_MODE `i_axi_a2x_2_A2X_BRESP_MODE
`endif 

`ifdef i_axi_a2x_2_A2X_BRESP_ORDER
  `define A2X_BRESP_ORDER `i_axi_a2x_2_A2X_BRESP_ORDER
`endif 

`ifdef i_axi_a2x_2_A2X_OSW_EN
  `define A2X_OSW_EN `i_axi_a2x_2_A2X_OSW_EN
`endif 

`ifdef i_axi_a2x_2_A2X_NUM_UWID
  `define A2X_NUM_UWID `i_axi_a2x_2_A2X_NUM_UWID
`endif 

`ifdef i_axi_a2x_2_A2X_SP_OSAW_LIMIT_P1
  `define A2X_SP_OSAW_LIMIT_P1 `i_axi_a2x_2_A2X_SP_OSAW_LIMIT_P1
`endif 

`ifdef i_axi_a2x_2_A2X_SP_OSAW_LIMIT
  `define A2X_SP_OSAW_LIMIT `i_axi_a2x_2_A2X_SP_OSAW_LIMIT
`endif 

`ifdef i_axi_a2x_2_A2X_OSAW_LIMIT
  `define A2X_OSAW_LIMIT `i_axi_a2x_2_A2X_OSAW_LIMIT
`endif 

`ifdef i_axi_a2x_2_A2X_PP_OSAW_LIMIT_P1
  `define A2X_PP_OSAW_LIMIT_P1 `i_axi_a2x_2_A2X_PP_OSAW_LIMIT_P1
`endif 

`ifdef i_axi_a2x_2_A2X_PP_OSAW_LIMIT
  `define A2X_PP_OSAW_LIMIT `i_axi_a2x_2_A2X_PP_OSAW_LIMIT
`endif 

`ifdef i_axi_a2x_2_A2X_B_OSW_LIMIT_P1
  `define A2X_B_OSW_LIMIT_P1 `i_axi_a2x_2_A2X_B_OSW_LIMIT_P1
`endif 

`ifdef i_axi_a2x_2_A2X_B_OSW_LIMIT
  `define A2X_B_OSW_LIMIT `i_axi_a2x_2_A2X_B_OSW_LIMIT
`endif 

`ifdef i_axi_a2x_2_A2X_OSW_LIMIT
  `define A2X_OSW_LIMIT `i_axi_a2x_2_A2X_OSW_LIMIT
`endif 

`ifdef i_axi_a2x_2_A2X_RBUF_MODE
  `define A2X_RBUF_MODE `i_axi_a2x_2_A2X_RBUF_MODE
`endif 

`ifdef i_axi_a2x_2_A2X_HCSNF_RLEN
  `define A2X_HCSNF_RLEN `i_axi_a2x_2_A2X_HCSNF_RLEN
`endif 

`ifdef i_axi_a2x_2_A2X_SNF_ARLEN_DFLT
  `define A2X_SNF_ARLEN_DFLT `i_axi_a2x_2_A2X_SNF_ARLEN_DFLT
`endif 

`ifdef i_axi_a2x_2_A2X_SNF_ARLEN_MIN
  `define A2X_SNF_ARLEN_MIN `i_axi_a2x_2_A2X_SNF_ARLEN_MIN
`endif 

`ifdef i_axi_a2x_2_A2X_AHB_RRECALL_DEPTH
  `define A2X_AHB_RRECALL_DEPTH `i_axi_a2x_2_A2X_AHB_RRECALL_DEPTH
`endif 

`ifdef i_axi_a2x_2_A2X_AHB_EBT_MODE
  `define A2X_AHB_EBT_MODE `i_axi_a2x_2_A2X_AHB_EBT_MODE
`endif 

`ifdef i_axi_a2x_2_A2X_HINCR_RBCNT_MIN
  `define A2X_HINCR_RBCNT_MIN `i_axi_a2x_2_A2X_HINCR_RBCNT_MIN
`endif 

`ifdef i_axi_a2x_2_A2X_HINCR_RBCNT_MAX
  `define A2X_HINCR_RBCNT_MAX `i_axi_a2x_2_A2X_HINCR_RBCNT_MAX
`endif 

`ifdef i_axi_a2x_2_A2X_LKMODE_MAX_PREFETCH
  `define A2X_LKMODE_MAX_PREFETCH `i_axi_a2x_2_A2X_LKMODE_MAX_PREFETCH
`endif 

`ifdef i_axi_a2x_2_A2X_HINCR_ARLEN_DFLT
  `define A2X_HINCR_ARLEN_DFLT `i_axi_a2x_2_A2X_HINCR_ARLEN_DFLT
`endif 

`ifdef i_axi_a2x_2_A2X_HINCR_ARLEN_MIN
  `define A2X_HINCR_ARLEN_MIN `i_axi_a2x_2_A2X_HINCR_ARLEN_MIN
`endif 

`ifdef i_axi_a2x_2_A2X_READ_INTLEV
  `define A2X_READ_INTLEV `i_axi_a2x_2_A2X_READ_INTLEV
`endif 

`ifdef i_axi_a2x_2_A2X_READ_ORDER
  `define A2X_READ_ORDER `i_axi_a2x_2_A2X_READ_ORDER
`endif 

`ifdef i_axi_a2x_2_SIM_REORDER
  `define SIM_REORDER `i_axi_a2x_2_SIM_REORDER
`endif 

`ifdef i_axi_a2x_2_A2X_OSR_EN
  `define A2X_OSR_EN `i_axi_a2x_2_A2X_OSR_EN
`endif 

`ifdef i_axi_a2x_2_A2X_NUM_URID
  `define A2X_NUM_URID `i_axi_a2x_2_A2X_NUM_URID
`endif 

`ifdef i_axi_a2x_2_A2X_OSR_LIMIT_P1
  `define A2X_OSR_LIMIT_P1 `i_axi_a2x_2_A2X_OSR_LIMIT_P1
`endif 

`ifdef i_axi_a2x_2_A2X_OSR_LIMIT
  `define A2X_OSR_LIMIT `i_axi_a2x_2_A2X_OSR_LIMIT
`endif 

`ifdef i_axi_a2x_2_A2X_A_UBW
  `define A2X_A_UBW `i_axi_a2x_2_A2X_A_UBW
`endif 

`ifdef i_axi_a2x_2_A2X_USER_SIGNAL_XFER_MODE
  `define A2X_USER_SIGNAL_XFER_MODE `i_axi_a2x_2_A2X_USER_SIGNAL_XFER_MODE
`endif 

`ifdef i_axi_a2x_2_A2X_WUSER_BITS_PER_BYTE
  `define A2X_WUSER_BITS_PER_BYTE `i_axi_a2x_2_A2X_WUSER_BITS_PER_BYTE
`endif 

`ifdef i_axi_a2x_2_A2X_RUSER_BITS_PER_BYTE
  `define A2X_RUSER_BITS_PER_BYTE `i_axi_a2x_2_A2X_RUSER_BITS_PER_BYTE
`endif 

`ifdef i_axi_a2x_2_A2X_W_UBW
  `define A2X_W_UBW `i_axi_a2x_2_A2X_W_UBW
`endif 

`ifdef i_axi_a2x_2_A2X_R_UBW
  `define A2X_R_UBW `i_axi_a2x_2_A2X_R_UBW
`endif 

`ifdef i_axi_a2x_2_A2X_AWSBW
  `define A2X_AWSBW `i_axi_a2x_2_A2X_AWSBW
`endif 

`ifdef i_axi_a2x_2_A2X_ARSBW
  `define A2X_ARSBW `i_axi_a2x_2_A2X_ARSBW
`endif 

`ifdef i_axi_a2x_2_A2X_WSBW
  `define A2X_WSBW `i_axi_a2x_2_A2X_WSBW
`endif 

`ifdef i_axi_a2x_2_A2X_RSBW
  `define A2X_RSBW `i_axi_a2x_2_A2X_RSBW
`endif 

`ifdef i_axi_a2x_2_A2X_BSBW
  `define A2X_BSBW `i_axi_a2x_2_A2X_BSBW
`endif 

`ifdef i_axi_a2x_2_A2X_INC_QOS
  `define A2X_INC_QOS `i_axi_a2x_2_A2X_INC_QOS
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_QOS
  `define A2X_HAS_QOS `i_axi_a2x_2_A2X_HAS_QOS
`endif 

`ifdef i_axi_a2x_2_A2X_INC_REGION
  `define A2X_INC_REGION `i_axi_a2x_2_A2X_INC_REGION
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_REGION
  `define A2X_HAS_REGION `i_axi_a2x_2_A2X_HAS_REGION
`endif 

`ifdef i_axi_a2x_2_A2X_AW_FIFO_DEPTH
  `define A2X_AW_FIFO_DEPTH `i_axi_a2x_2_A2X_AW_FIFO_DEPTH
`endif 

`ifdef i_axi_a2x_2_A2X_WD_FIFO_DEPTH
  `define A2X_WD_FIFO_DEPTH `i_axi_a2x_2_A2X_WD_FIFO_DEPTH
`endif 

`ifdef i_axi_a2x_2_A2X_BRESP_FIFO_DEPTH
  `define A2X_BRESP_FIFO_DEPTH `i_axi_a2x_2_A2X_BRESP_FIFO_DEPTH
`endif 

`ifdef i_axi_a2x_2_A2X_AR_FIFO_DEPTH
  `define A2X_AR_FIFO_DEPTH `i_axi_a2x_2_A2X_AR_FIFO_DEPTH
`endif 

`ifdef i_axi_a2x_2_A2X_RD_FIFO_DEPTH
  `define A2X_RD_FIFO_DEPTH `i_axi_a2x_2_A2X_RD_FIFO_DEPTH
`endif 

`ifdef i_axi_a2x_2_A2X_LK_RD_FIFO_DEPTH
  `define A2X_LK_RD_FIFO_DEPTH `i_axi_a2x_2_A2X_LK_RD_FIFO_DEPTH
`endif 

`ifdef i_axi_a2x_2_A2X_AUTO_LINK_SPLIT_MODE
  `define A2X_AUTO_LINK_SPLIT_MODE `i_axi_a2x_2_A2X_AUTO_LINK_SPLIT_MODE
`endif 

`ifdef i_axi_a2x_2_A2X_AR_SP_PIPELINE
  `define A2X_AR_SP_PIPELINE `i_axi_a2x_2_A2X_AR_SP_PIPELINE
`endif 

`ifdef i_axi_a2x_2_A2X_AW_SP_PIPELINE
  `define A2X_AW_SP_PIPELINE `i_axi_a2x_2_A2X_AW_SP_PIPELINE
`endif 

`ifdef i_axi_a2x_2_A2X_RS_AR_TMO
  `define A2X_RS_AR_TMO `i_axi_a2x_2_A2X_RS_AR_TMO
`endif 

`ifdef i_axi_a2x_2_A2X_RS_AW_TMO
  `define A2X_RS_AW_TMO `i_axi_a2x_2_A2X_RS_AW_TMO
`endif 

`ifdef i_axi_a2x_2_A2X_RS_R_TMO
  `define A2X_RS_R_TMO `i_axi_a2x_2_A2X_RS_R_TMO
`endif 

`ifdef i_axi_a2x_2_A2X_RS_W_TMO
  `define A2X_RS_W_TMO `i_axi_a2x_2_A2X_RS_W_TMO
`endif 

`ifdef i_axi_a2x_2_A2X_RS_B_TMO
  `define A2X_RS_B_TMO `i_axi_a2x_2_A2X_RS_B_TMO
`endif 

`ifdef i_axi_a2x_2_A2X_AHB_LOCKED
  `define A2X_AHB_LOCKED `i_axi_a2x_2_A2X_AHB_LOCKED
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_LOCKED
  `define A2X_HAS_LOCKED `i_axi_a2x_2_A2X_HAS_LOCKED
`endif 

`ifdef i_axi_a2x_2_A2X_INT_NUM_AHBM
  `define A2X_INT_NUM_AHBM `i_axi_a2x_2_A2X_INT_NUM_AHBM
`endif 

`ifdef i_axi_a2x_2_A2X_UPSIZE
  `define A2X_UPSIZE `i_axi_a2x_2_A2X_UPSIZE
`endif 

`ifdef i_axi_a2x_2_A2X_DOWNSIZE
  `define A2X_DOWNSIZE `i_axi_a2x_2_A2X_DOWNSIZE
`endif 

`ifdef i_axi_a2x_2_A2X_IS_UPSIZED
  `define A2X_IS_UPSIZED `i_axi_a2x_2_A2X_IS_UPSIZED
`endif 

`ifdef i_axi_a2x_2_A2X_IS_DOWNSIZED
  `define A2X_IS_DOWNSIZED `i_axi_a2x_2_A2X_IS_DOWNSIZED
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_RBUF
  `define A2X_HAS_RBUF `i_axi_a2x_2_A2X_HAS_RBUF
`endif 

`ifdef i_axi_a2x_2_A2X_IS_EQSIZED
  `define A2X_IS_EQSIZED `i_axi_a2x_2_A2X_IS_EQSIZED
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_NBUF_MODE
  `define A2X_HAS_NBUF_MODE `i_axi_a2x_2_A2X_HAS_NBUF_MODE
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_HINCR_HCBCNT
  `define A2X_HAS_HINCR_HCBCNT `i_axi_a2x_2_A2X_HAS_HINCR_HCBCNT
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_SINGLE_RBCNT
  `define A2X_HAS_SINGLE_RBCNT `i_axi_a2x_2_A2X_HAS_SINGLE_RBCNT
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_SINGLE_WBCNT
  `define A2X_HAS_SINGLE_WBCNT `i_axi_a2x_2_A2X_HAS_SINGLE_WBCNT
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_CNT_M1
  `define A2X_HAS_CNT_M1 `i_axi_a2x_2_A2X_HAS_CNT_M1
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_CNT_M2
  `define A2X_HAS_CNT_M2 `i_axi_a2x_2_A2X_HAS_CNT_M2
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_CNT_M3
  `define A2X_HAS_CNT_M3 `i_axi_a2x_2_A2X_HAS_CNT_M3
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_CNT_M4
  `define A2X_HAS_CNT_M4 `i_axi_a2x_2_A2X_HAS_CNT_M4
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_CNT_M5
  `define A2X_HAS_CNT_M5 `i_axi_a2x_2_A2X_HAS_CNT_M5
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_CNT_M6
  `define A2X_HAS_CNT_M6 `i_axi_a2x_2_A2X_HAS_CNT_M6
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_CNT_M7
  `define A2X_HAS_CNT_M7 `i_axi_a2x_2_A2X_HAS_CNT_M7
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_CNT_M8
  `define A2X_HAS_CNT_M8 `i_axi_a2x_2_A2X_HAS_CNT_M8
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_CNT_M9
  `define A2X_HAS_CNT_M9 `i_axi_a2x_2_A2X_HAS_CNT_M9
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_CNT_M10
  `define A2X_HAS_CNT_M10 `i_axi_a2x_2_A2X_HAS_CNT_M10
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_CNT_M11
  `define A2X_HAS_CNT_M11 `i_axi_a2x_2_A2X_HAS_CNT_M11
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_CNT_M12
  `define A2X_HAS_CNT_M12 `i_axi_a2x_2_A2X_HAS_CNT_M12
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_CNT_M13
  `define A2X_HAS_CNT_M13 `i_axi_a2x_2_A2X_HAS_CNT_M13
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_CNT_M14
  `define A2X_HAS_CNT_M14 `i_axi_a2x_2_A2X_HAS_CNT_M14
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_CNT_M15
  `define A2X_HAS_CNT_M15 `i_axi_a2x_2_A2X_HAS_CNT_M15
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_LOWPWR_IF
  `define A2X_HAS_LOWPWR_IF `i_axi_a2x_2_A2X_HAS_LOWPWR_IF
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_USER_SIGNAL_XFER_MODE
  `define A2X_HAS_USER_SIGNAL_XFER_MODE `i_axi_a2x_2_A2X_HAS_USER_SIGNAL_XFER_MODE
`endif 

`ifdef i_axi_a2x_2_A2X_INT_HASBW
  `define A2X_INT_HASBW `i_axi_a2x_2_A2X_INT_HASBW
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_HASB
  `define A2X_HAS_HASB `i_axi_a2x_2_A2X_HAS_HASB
`endif 

`ifdef i_axi_a2x_2_A2X_INT_HWSBW
  `define A2X_INT_HWSBW `i_axi_a2x_2_A2X_INT_HWSBW
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_HWSB
  `define A2X_HAS_HWSB `i_axi_a2x_2_A2X_HAS_HWSB
`endif 

`ifdef i_axi_a2x_2_A2X_INT_HRSBW
  `define A2X_INT_HRSBW `i_axi_a2x_2_A2X_INT_HRSBW
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_HRSB
  `define A2X_HAS_HRSB `i_axi_a2x_2_A2X_HAS_HRSB
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_AWSB
  `define A2X_HAS_AWSB `i_axi_a2x_2_A2X_HAS_AWSB
`endif 

`ifdef i_axi_a2x_2_A2X_INT_AWSBW
  `define A2X_INT_AWSBW `i_axi_a2x_2_A2X_INT_AWSBW
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_WSB
  `define A2X_HAS_WSB `i_axi_a2x_2_A2X_HAS_WSB
`endif 

`ifdef i_axi_a2x_2_A2X_INT_WSBW
  `define A2X_INT_WSBW `i_axi_a2x_2_A2X_INT_WSBW
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_ARSB
  `define A2X_HAS_ARSB `i_axi_a2x_2_A2X_HAS_ARSB
`endif 

`ifdef i_axi_a2x_2_A2X_INT_ARSBW
  `define A2X_INT_ARSBW `i_axi_a2x_2_A2X_INT_ARSBW
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_RSB
  `define A2X_HAS_RSB `i_axi_a2x_2_A2X_HAS_RSB
`endif 

`ifdef i_axi_a2x_2_A2X_INT_RSBW
  `define A2X_INT_RSBW `i_axi_a2x_2_A2X_INT_RSBW
`endif 

`ifdef i_axi_a2x_2_A2X_HAS_BSB
  `define A2X_HAS_BSB `i_axi_a2x_2_A2X_HAS_BSB
`endif 

`ifdef i_axi_a2x_2_A2X_INT_BSBW
  `define A2X_INT_BSBW `i_axi_a2x_2_A2X_INT_BSBW
`endif 

`ifdef i_axi_a2x_2_A2X_PP_IS_AHB
  `define A2X_PP_IS_AHB `i_axi_a2x_2_A2X_PP_IS_AHB
`endif 

`ifdef i_axi_a2x_2_A2X_PP_IS_AXI
  `define A2X_PP_IS_AXI `i_axi_a2x_2_A2X_PP_IS_AXI
`endif 

`ifdef i_axi_a2x_2_A2X_CLK_IS_SYNC
  `define A2X_CLK_IS_SYNC `i_axi_a2x_2_A2X_CLK_IS_SYNC
`endif 

`ifdef i_axi_a2x_2_A2X_AW_FIFO_DEPTH_LOG2
  `define A2X_AW_FIFO_DEPTH_LOG2 `i_axi_a2x_2_A2X_AW_FIFO_DEPTH_LOG2
`endif 

`ifdef i_axi_a2x_2_A2X_AR_FIFO_DEPTH_LOG2
  `define A2X_AR_FIFO_DEPTH_LOG2 `i_axi_a2x_2_A2X_AR_FIFO_DEPTH_LOG2
`endif 

`ifdef i_axi_a2x_2_A2X_BRESP_FIFO_DEPTH_LOG2
  `define A2X_BRESP_FIFO_DEPTH_LOG2 `i_axi_a2x_2_A2X_BRESP_FIFO_DEPTH_LOG2
`endif 

`ifdef i_axi_a2x_2_A2X_WD_FIFO_DEPTH_LOG2
  `define A2X_WD_FIFO_DEPTH_LOG2 `i_axi_a2x_2_A2X_WD_FIFO_DEPTH_LOG2
`endif 

`ifdef i_axi_a2x_2_A2X_RD_FIFO_DEPTH_LOG2
  `define A2X_RD_FIFO_DEPTH_LOG2 `i_axi_a2x_2_A2X_RD_FIFO_DEPTH_LOG2
`endif 

`ifdef i_axi_a2x_2_A2X_B_OSW_LIMIT_LOG2
  `define A2X_B_OSW_LIMIT_LOG2 `i_axi_a2x_2_A2X_B_OSW_LIMIT_LOG2
`endif 

`ifdef i_axi_a2x_2_A2X_PP_OSAW_LIMIT_LOG2
  `define A2X_PP_OSAW_LIMIT_LOG2 `i_axi_a2x_2_A2X_PP_OSAW_LIMIT_LOG2
`endif 

`ifdef i_axi_a2x_2_A2X_SP_OSAW_LIMIT_LOG2
  `define A2X_SP_OSAW_LIMIT_LOG2 `i_axi_a2x_2_A2X_SP_OSAW_LIMIT_LOG2
`endif 

`ifdef i_axi_a2x_2_A2X_OSR_LIMIT_LOG2
  `define A2X_OSR_LIMIT_LOG2 `i_axi_a2x_2_A2X_OSR_LIMIT_LOG2
`endif 

`ifdef i_axi_a2x_2_A2X_LK_RD_FIFO_DEPTH_LOG2
  `define A2X_LK_RD_FIFO_DEPTH_LOG2 `i_axi_a2x_2_A2X_LK_RD_FIFO_DEPTH_LOG2
`endif 

`ifdef i_axi_a2x_2_A2X_PP_DW_LOG2
  `define A2X_PP_DW_LOG2 `i_axi_a2x_2_A2X_PP_DW_LOG2
`endif 

`ifdef i_axi_a2x_2_A2X_SP_DW_LOG2
  `define A2X_SP_DW_LOG2 `i_axi_a2x_2_A2X_SP_DW_LOG2
`endif 

`ifdef i_axi_a2x_2_A2X_PP_NUM_BYTES
  `define A2X_PP_NUM_BYTES `i_axi_a2x_2_A2X_PP_NUM_BYTES
`endif 

`ifdef i_axi_a2x_2_A2X_PP_WSTRB_DW
  `define A2X_PP_WSTRB_DW `i_axi_a2x_2_A2X_PP_WSTRB_DW
`endif 

`ifdef i_axi_a2x_2_A2X_SP_NUM_BYTES
  `define A2X_SP_NUM_BYTES `i_axi_a2x_2_A2X_SP_NUM_BYTES
`endif 

`ifdef i_axi_a2x_2_A2X_SP_WSTRB_DW
  `define A2X_SP_WSTRB_DW `i_axi_a2x_2_A2X_SP_WSTRB_DW
`endif 

`ifdef i_axi_a2x_2_A2X_PP_MAX_SIZE
  `define A2X_PP_MAX_SIZE `i_axi_a2x_2_A2X_PP_MAX_SIZE
`endif 

`ifdef i_axi_a2x_2_A2X_SP_MAX_SIZE
  `define A2X_SP_MAX_SIZE `i_axi_a2x_2_A2X_SP_MAX_SIZE
`endif 

`ifdef i_axi_a2x_2_A2X_MAX_PP_TOTAL_BYTES
  `define A2X_MAX_PP_TOTAL_BYTES `i_axi_a2x_2_A2X_MAX_PP_TOTAL_BYTES
`endif 

`ifdef i_axi_a2x_2_A2X_MAX_SP_TOTAL_BYTES
  `define A2X_MAX_SP_TOTAL_BYTES `i_axi_a2x_2_A2X_MAX_SP_TOTAL_BYTES
`endif 

`ifdef i_axi_a2x_2_A2X_MAX_TOTAL_BYTES
  `define A2X_MAX_TOTAL_BYTES `i_axi_a2x_2_A2X_MAX_TOTAL_BYTES
`endif 

`ifdef i_axi_a2x_2_A2X_MAX_TOTAL_BYTES_LOG2
  `define A2X_MAX_TOTAL_BYTES_LOG2 `i_axi_a2x_2_A2X_MAX_TOTAL_BYTES_LOG2
`endif 

`ifdef i_axi_a2x_2_A2X_PP_NUM_BYTES_LOG2
  `define A2X_PP_NUM_BYTES_LOG2 `i_axi_a2x_2_A2X_PP_NUM_BYTES_LOG2
`endif 

`ifdef i_axi_a2x_2_A2X_SP_NUM_BYTES_LOG2
  `define A2X_SP_NUM_BYTES_LOG2 `i_axi_a2x_2_A2X_SP_NUM_BYTES_LOG2
`endif 

`ifdef i_axi_a2x_2_A2X_PP_DW_16
  `define A2X_PP_DW_16 `i_axi_a2x_2_A2X_PP_DW_16
`endif 

`ifdef i_axi_a2x_2_A2X_PP_DW_32
  `define A2X_PP_DW_32 `i_axi_a2x_2_A2X_PP_DW_32
`endif 

`ifdef i_axi_a2x_2_A2X_PP_DW_64
  `define A2X_PP_DW_64 `i_axi_a2x_2_A2X_PP_DW_64
`endif 

`ifdef i_axi_a2x_2_A2X_PP_DW_128
  `define A2X_PP_DW_128 `i_axi_a2x_2_A2X_PP_DW_128
`endif 

`ifdef i_axi_a2x_2_A2X_PP_DW_256
  `define A2X_PP_DW_256 `i_axi_a2x_2_A2X_PP_DW_256
`endif 

`ifdef i_axi_a2x_2_A2X_PP_DW_512
  `define A2X_PP_DW_512 `i_axi_a2x_2_A2X_PP_DW_512
`endif 

`ifdef i_axi_a2x_2_A2X_PP_DW_1024
  `define A2X_PP_DW_1024 `i_axi_a2x_2_A2X_PP_DW_1024
`endif 

`ifdef i_axi_a2x_2_A2X_SP_DW_32
  `define A2X_SP_DW_32 `i_axi_a2x_2_A2X_SP_DW_32
`endif 

`ifdef i_axi_a2x_2_A2X_SP_DW_64
  `define A2X_SP_DW_64 `i_axi_a2x_2_A2X_SP_DW_64
`endif 

`ifdef i_axi_a2x_2_A2X_SP_DW_128
  `define A2X_SP_DW_128 `i_axi_a2x_2_A2X_SP_DW_128
`endif 

`ifdef i_axi_a2x_2_A2X_SP_DW_256
  `define A2X_SP_DW_256 `i_axi_a2x_2_A2X_SP_DW_256
`endif 

`ifdef i_axi_a2x_2_A2X_SP_DW_512
  `define A2X_SP_DW_512 `i_axi_a2x_2_A2X_SP_DW_512
`endif 

`ifdef i_axi_a2x_2_A2X_SP_DW_1024
  `define A2X_SP_DW_1024 `i_axi_a2x_2_A2X_SP_DW_1024
`endif 

`ifdef i_axi_a2x_2_A2X_DS_RATIO_2
  `define A2X_DS_RATIO_2 `i_axi_a2x_2_A2X_DS_RATIO_2
`endif 

`ifdef i_axi_a2x_2_A2X_DS_RATIO_4
  `define A2X_DS_RATIO_4 `i_axi_a2x_2_A2X_DS_RATIO_4
`endif 

`ifdef i_axi_a2x_2_A2X_DS_RATIO_8
  `define A2X_DS_RATIO_8 `i_axi_a2x_2_A2X_DS_RATIO_8
`endif 

`ifdef i_axi_a2x_2_DWC_NO_TST_MODE
  `define DWC_NO_TST_MODE `i_axi_a2x_2_DWC_NO_TST_MODE
`endif 

`ifdef i_axi_a2x_2_DWC_NO_CDC_INIT
  `define DWC_NO_CDC_INIT `i_axi_a2x_2_DWC_NO_CDC_INIT
`endif 

`ifdef i_axi_a2x_2_A2X_SIM_SEED
  `define A2X_SIM_SEED `i_axi_a2x_2_A2X_SIM_SEED
`endif 

`ifdef i_axi_a2x_2_A2X_SIM_APB_CLK_PERIOD
  `define A2X_SIM_APB_CLK_PERIOD `i_axi_a2x_2_A2X_SIM_APB_CLK_PERIOD
`endif 

`ifdef i_axi_a2x_2_A2X_SIM_PP_CLK_PERIOD
  `define A2X_SIM_PP_CLK_PERIOD `i_axi_a2x_2_A2X_SIM_PP_CLK_PERIOD
`endif 

`ifdef i_axi_a2x_2_A2X_SIM_SP_CLK_PERIOD
  `define A2X_SIM_SP_CLK_PERIOD `i_axi_a2x_2_A2X_SIM_SP_CLK_PERIOD
`endif 

`ifdef i_axi_a2x_2_A2X_SP_CLK_SKEW
  `define A2X_SP_CLK_SKEW `i_axi_a2x_2_A2X_SP_CLK_SKEW
`endif 

`ifdef i_axi_a2x_2_A2X_INACTIVE_VAL
  `define A2X_INACTIVE_VAL `i_axi_a2x_2_A2X_INACTIVE_VAL
`endif 

`ifdef i_axi_a2x_2_A2X_ASYNC_CLKS
  `define A2X_ASYNC_CLKS `i_axi_a2x_2_A2X_ASYNC_CLKS
`endif 

`ifdef i_axi_a2x_2_A2X_DUAL_CLK
  `define A2X_DUAL_CLK `i_axi_a2x_2_A2X_DUAL_CLK
`endif 

`ifdef i_axi_a2x_2_A2X_N_TESTCASE_DUPLICATION
  `define A2X_N_TESTCASE_DUPLICATION `i_axi_a2x_2_A2X_N_TESTCASE_DUPLICATION
`endif 

`ifdef i_axi_a2x_2_A2X_PRIMEPOWER_SIM
  `define A2X_PRIMEPOWER_SIM `i_axi_a2x_2_A2X_PRIMEPOWER_SIM
`endif 

`ifdef i_axi_a2x_2_A2X_SIM_IS_PRIMEPOWER
  `define A2X_SIM_IS_PRIMEPOWER `i_axi_a2x_2_A2X_SIM_IS_PRIMEPOWER
`endif 

`ifdef i_axi_a2x_2_A2X_VERIF_EN
  `define A2X_VERIF_EN `i_axi_a2x_2_A2X_VERIF_EN
`endif 

`ifdef i_axi_a2x_2_A2X_HRESPW
  `define A2X_HRESPW `i_axi_a2x_2_A2X_HRESPW
`endif 

`ifdef i_axi_a2x_2_A2X_HRESP_WIDTH_2
  `define A2X_HRESP_WIDTH_2 `i_axi_a2x_2_A2X_HRESP_WIDTH_2
`endif 

`ifdef i_axi_a2x_2___GUARD__DW_AXI_A2X_BCM_PARAMS__VH__
  `define __GUARD__DW_AXI_A2X_BCM_PARAMS__VH__ `i_axi_a2x_2___GUARD__DW_AXI_A2X_BCM_PARAMS__VH__
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM00_AND
  `define DW_AXI_A2X_RM_BCM00_AND `i_axi_a2x_2_DW_AXI_A2X_RM_BCM00_AND
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM00_ATPG_MX
  `define DW_AXI_A2X_RM_BCM00_ATPG_MX `i_axi_a2x_2_DW_AXI_A2X_RM_BCM00_ATPG_MX
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM00_CK_AND
  `define DW_AXI_A2X_RM_BCM00_CK_AND `i_axi_a2x_2_DW_AXI_A2X_RM_BCM00_CK_AND
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM00_CK_BUF
  `define DW_AXI_A2X_RM_BCM00_CK_BUF `i_axi_a2x_2_DW_AXI_A2X_RM_BCM00_CK_BUF
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM00_CK_GT_LAT
  `define DW_AXI_A2X_RM_BCM00_CK_GT_LAT `i_axi_a2x_2_DW_AXI_A2X_RM_BCM00_CK_GT_LAT
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM00_CK_MX
  `define DW_AXI_A2X_RM_BCM00_CK_MX `i_axi_a2x_2_DW_AXI_A2X_RM_BCM00_CK_MX
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM00_CK_OR
  `define DW_AXI_A2X_RM_BCM00_CK_OR `i_axi_a2x_2_DW_AXI_A2X_RM_BCM00_CK_OR
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM00_MAJ
  `define DW_AXI_A2X_RM_BCM00_MAJ `i_axi_a2x_2_DW_AXI_A2X_RM_BCM00_MAJ
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM00_MX
  `define DW_AXI_A2X_RM_BCM00_MX `i_axi_a2x_2_DW_AXI_A2X_RM_BCM00_MX
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM00_OR
  `define DW_AXI_A2X_RM_BCM00_OR `i_axi_a2x_2_DW_AXI_A2X_RM_BCM00_OR
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM01
  `define DW_AXI_A2X_RM_BCM01 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM01
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM02
  `define DW_AXI_A2X_RM_BCM02 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM02
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM03
  `define DW_AXI_A2X_RM_BCM03 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM03
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM04
  `define DW_AXI_A2X_RM_BCM04 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM04
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM05
  `define DW_AXI_A2X_RM_BCM05 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM05
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM05_ATV
  `define DW_AXI_A2X_RM_BCM05_ATV `i_axi_a2x_2_DW_AXI_A2X_RM_BCM05_ATV
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM05_CF
  `define DW_AXI_A2X_RM_BCM05_CF `i_axi_a2x_2_DW_AXI_A2X_RM_BCM05_CF
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM05_EF
  `define DW_AXI_A2X_RM_BCM05_EF `i_axi_a2x_2_DW_AXI_A2X_RM_BCM05_EF
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM05_EF_ATV
  `define DW_AXI_A2X_RM_BCM05_EF_ATV `i_axi_a2x_2_DW_AXI_A2X_RM_BCM05_EF_ATV
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM06
  `define DW_AXI_A2X_RM_BCM06 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM06
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM06_ATV
  `define DW_AXI_A2X_RM_BCM06_ATV `i_axi_a2x_2_DW_AXI_A2X_RM_BCM06_ATV
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM07
  `define DW_AXI_A2X_RM_BCM07 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM07
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM07_ATV
  `define DW_AXI_A2X_RM_BCM07_ATV `i_axi_a2x_2_DW_AXI_A2X_RM_BCM07_ATV
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM07_EF
  `define DW_AXI_A2X_RM_BCM07_EF `i_axi_a2x_2_DW_AXI_A2X_RM_BCM07_EF
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM07_EF_ATV
  `define DW_AXI_A2X_RM_BCM07_EF_ATV `i_axi_a2x_2_DW_AXI_A2X_RM_BCM07_EF_ATV
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM07_EFES
  `define DW_AXI_A2X_RM_BCM07_EFES `i_axi_a2x_2_DW_AXI_A2X_RM_BCM07_EFES
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM07_RS
  `define DW_AXI_A2X_RM_BCM07_RS `i_axi_a2x_2_DW_AXI_A2X_RM_BCM07_RS
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM08
  `define DW_AXI_A2X_RM_BCM08 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM08
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM09
  `define DW_AXI_A2X_RM_BCM09 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM09
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM09_DP
  `define DW_AXI_A2X_RM_BCM09_DP `i_axi_a2x_2_DW_AXI_A2X_RM_BCM09_DP
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM09_ECC
  `define DW_AXI_A2X_RM_BCM09_ECC `i_axi_a2x_2_DW_AXI_A2X_RM_BCM09_ECC
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM10
  `define DW_AXI_A2X_RM_BCM10 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM10
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM11
  `define DW_AXI_A2X_RM_BCM11 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM11
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM12
  `define DW_AXI_A2X_RM_BCM12 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM12
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM14
  `define DW_AXI_A2X_RM_BCM14 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM14
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM15
  `define DW_AXI_A2X_RM_BCM15 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM15
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM16
  `define DW_AXI_A2X_RM_BCM16 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM16
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM17
  `define DW_AXI_A2X_RM_BCM17 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM17
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM18_GEN
  `define DW_AXI_A2X_RM_BCM18_GEN `i_axi_a2x_2_DW_AXI_A2X_RM_BCM18_GEN
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM18_MON
  `define DW_AXI_A2X_RM_BCM18_MON `i_axi_a2x_2_DW_AXI_A2X_RM_BCM18_MON
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM18_PGEN
  `define DW_AXI_A2X_RM_BCM18_PGEN `i_axi_a2x_2_DW_AXI_A2X_RM_BCM18_PGEN
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM18_PGENA
  `define DW_AXI_A2X_RM_BCM18_PGENA `i_axi_a2x_2_DW_AXI_A2X_RM_BCM18_PGENA
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM18_PMON
  `define DW_AXI_A2X_RM_BCM18_PMON `i_axi_a2x_2_DW_AXI_A2X_RM_BCM18_PMON
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM18_RS
  `define DW_AXI_A2X_RM_BCM18_RS `i_axi_a2x_2_DW_AXI_A2X_RM_BCM18_RS
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM19_INTR
  `define DW_AXI_A2X_RM_BCM19_INTR `i_axi_a2x_2_DW_AXI_A2X_RM_BCM19_INTR
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM19_TRGT
  `define DW_AXI_A2X_RM_BCM19_TRGT `i_axi_a2x_2_DW_AXI_A2X_RM_BCM19_TRGT
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM21
  `define DW_AXI_A2X_RM_BCM21 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM21
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM21_ATV
  `define DW_AXI_A2X_RM_BCM21_ATV `i_axi_a2x_2_DW_AXI_A2X_RM_BCM21_ATV
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM21_NEO
  `define DW_AXI_A2X_RM_BCM21_NEO `i_axi_a2x_2_DW_AXI_A2X_RM_BCM21_NEO
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM21_TGL
  `define DW_AXI_A2X_RM_BCM21_TGL `i_axi_a2x_2_DW_AXI_A2X_RM_BCM21_TGL
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM22
  `define DW_AXI_A2X_RM_BCM22 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM22
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM22_ATV
  `define DW_AXI_A2X_RM_BCM22_ATV `i_axi_a2x_2_DW_AXI_A2X_RM_BCM22_ATV
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM23
  `define DW_AXI_A2X_RM_BCM23 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM23
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM23_ATV
  `define DW_AXI_A2X_RM_BCM23_ATV `i_axi_a2x_2_DW_AXI_A2X_RM_BCM23_ATV
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM23_C
  `define DW_AXI_A2X_RM_BCM23_C `i_axi_a2x_2_DW_AXI_A2X_RM_BCM23_C
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM24
  `define DW_AXI_A2X_RM_BCM24 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM24
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM24_AP
  `define DW_AXI_A2X_RM_BCM24_AP `i_axi_a2x_2_DW_AXI_A2X_RM_BCM24_AP
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM25
  `define DW_AXI_A2X_RM_BCM25 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM25
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM25_ATV
  `define DW_AXI_A2X_RM_BCM25_ATV `i_axi_a2x_2_DW_AXI_A2X_RM_BCM25_ATV
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM25_C
  `define DW_AXI_A2X_RM_BCM25_C `i_axi_a2x_2_DW_AXI_A2X_RM_BCM25_C
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM26
  `define DW_AXI_A2X_RM_BCM26 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM26
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM26_ATV
  `define DW_AXI_A2X_RM_BCM26_ATV `i_axi_a2x_2_DW_AXI_A2X_RM_BCM26_ATV
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM27
  `define DW_AXI_A2X_RM_BCM27 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM27
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM28
  `define DW_AXI_A2X_RM_BCM28 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM28
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM29
  `define DW_AXI_A2X_RM_BCM29 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM29
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM31_P2D_FIFOMEM
  `define DW_AXI_A2X_RM_BCM31_P2D_FIFOMEM `i_axi_a2x_2_DW_AXI_A2X_RM_BCM31_P2D_FIFOMEM
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM31_P2D_RD
  `define DW_AXI_A2X_RM_BCM31_P2D_RD `i_axi_a2x_2_DW_AXI_A2X_RM_BCM31_P2D_RD
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM31_P2D_WR
  `define DW_AXI_A2X_RM_BCM31_P2D_WR `i_axi_a2x_2_DW_AXI_A2X_RM_BCM31_P2D_WR
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM32_A
  `define DW_AXI_A2X_RM_BCM32_A `i_axi_a2x_2_DW_AXI_A2X_RM_BCM32_A
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM32_C
  `define DW_AXI_A2X_RM_BCM32_C `i_axi_a2x_2_DW_AXI_A2X_RM_BCM32_C
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM33_63_7_64_0
  `define DW_AXI_A2X_RM_BCM33_63_7_64_0 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM33_63_7_64_0
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM35
  `define DW_AXI_A2X_RM_BCM35 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM35
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM35_T
  `define DW_AXI_A2X_RM_BCM35_T `i_axi_a2x_2_DW_AXI_A2X_RM_BCM35_T
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM36
  `define DW_AXI_A2X_RM_BCM36 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM36
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM36_ACK
  `define DW_AXI_A2X_RM_BCM36_ACK `i_axi_a2x_2_DW_AXI_A2X_RM_BCM36_ACK
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM36_NHS
  `define DW_AXI_A2X_RM_BCM36_NHS `i_axi_a2x_2_DW_AXI_A2X_RM_BCM36_NHS
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM36_TGL
  `define DW_AXI_A2X_RM_BCM36_TGL `i_axi_a2x_2_DW_AXI_A2X_RM_BCM36_TGL
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM36_TGL_DO
  `define DW_AXI_A2X_RM_BCM36_TGL_DO `i_axi_a2x_2_DW_AXI_A2X_RM_BCM36_TGL_DO
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM36_TGL_PLS
  `define DW_AXI_A2X_RM_BCM36_TGL_PLS `i_axi_a2x_2_DW_AXI_A2X_RM_BCM36_TGL_PLS
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM36_TGL_PLS_DO
  `define DW_AXI_A2X_RM_BCM36_TGL_PLS_DO `i_axi_a2x_2_DW_AXI_A2X_RM_BCM36_TGL_PLS_DO
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM37
  `define DW_AXI_A2X_RM_BCM37 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM37
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM38
  `define DW_AXI_A2X_RM_BCM38 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM38
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM38_ADP
  `define DW_AXI_A2X_RM_BCM38_ADP `i_axi_a2x_2_DW_AXI_A2X_RM_BCM38_ADP
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM38_AP
  `define DW_AXI_A2X_RM_BCM38_AP `i_axi_a2x_2_DW_AXI_A2X_RM_BCM38_AP
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM38_ECC
  `define DW_AXI_A2X_RM_BCM38_ECC `i_axi_a2x_2_DW_AXI_A2X_RM_BCM38_ECC
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM39
  `define DW_AXI_A2X_RM_BCM39 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM39
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM40
  `define DW_AXI_A2X_RM_BCM40 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM40
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM41
  `define DW_AXI_A2X_RM_BCM41 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM41
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM41_NEO
  `define DW_AXI_A2X_RM_BCM41_NEO `i_axi_a2x_2_DW_AXI_A2X_RM_BCM41_NEO
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM43
  `define DW_AXI_A2X_RM_BCM43 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM43
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM43_NRO
  `define DW_AXI_A2X_RM_BCM43_NRO `i_axi_a2x_2_DW_AXI_A2X_RM_BCM43_NRO
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM44
  `define DW_AXI_A2X_RM_BCM44 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM44
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM44_NRO
  `define DW_AXI_A2X_RM_BCM44_NRO `i_axi_a2x_2_DW_AXI_A2X_RM_BCM44_NRO
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_GN_D_A
  `define DW_AXI_A2X_RM_BCM45_GN_D_A `i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_GN_D_A
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_GN_D_AA
  `define DW_AXI_A2X_RM_BCM45_GN_D_AA `i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_GN_D_AA
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_GN_D_B
  `define DW_AXI_A2X_RM_BCM45_GN_D_B `i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_GN_D_B
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_GN_D_C
  `define DW_AXI_A2X_RM_BCM45_GN_D_C `i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_GN_D_C
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_GN_D_D
  `define DW_AXI_A2X_RM_BCM45_GN_D_D `i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_GN_D_D
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_GN_D_E
  `define DW_AXI_A2X_RM_BCM45_GN_D_E `i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_GN_D_E
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_GN_D_F
  `define DW_AXI_A2X_RM_BCM45_GN_D_F `i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_GN_D_F
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_MN_D_A
  `define DW_AXI_A2X_RM_BCM45_MN_D_A `i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_MN_D_A
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_MN_D_AA
  `define DW_AXI_A2X_RM_BCM45_MN_D_AA `i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_MN_D_AA
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_MN_D_B
  `define DW_AXI_A2X_RM_BCM45_MN_D_B `i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_MN_D_B
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_MN_D_C
  `define DW_AXI_A2X_RM_BCM45_MN_D_C `i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_MN_D_C
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_MN_D_D
  `define DW_AXI_A2X_RM_BCM45_MN_D_D `i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_MN_D_D
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_MN_D_E
  `define DW_AXI_A2X_RM_BCM45_MN_D_E `i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_MN_D_E
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_MN_D_F
  `define DW_AXI_A2X_RM_BCM45_MN_D_F `i_axi_a2x_2_DW_AXI_A2X_RM_BCM45_MN_D_F
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM46_A
  `define DW_AXI_A2X_RM_BCM46_A `i_axi_a2x_2_DW_AXI_A2X_RM_BCM46_A
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM46_AA
  `define DW_AXI_A2X_RM_BCM46_AA `i_axi_a2x_2_DW_AXI_A2X_RM_BCM46_AA
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM46_B
  `define DW_AXI_A2X_RM_BCM46_B `i_axi_a2x_2_DW_AXI_A2X_RM_BCM46_B
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM46_B_32A
  `define DW_AXI_A2X_RM_BCM46_B_32A `i_axi_a2x_2_DW_AXI_A2X_RM_BCM46_B_32A
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM46_C
  `define DW_AXI_A2X_RM_BCM46_C `i_axi_a2x_2_DW_AXI_A2X_RM_BCM46_C
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM46_C_64A
  `define DW_AXI_A2X_RM_BCM46_C_64A `i_axi_a2x_2_DW_AXI_A2X_RM_BCM46_C_64A
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM46_D
  `define DW_AXI_A2X_RM_BCM46_D `i_axi_a2x_2_DW_AXI_A2X_RM_BCM46_D
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM46_D_128A
  `define DW_AXI_A2X_RM_BCM46_D_128A `i_axi_a2x_2_DW_AXI_A2X_RM_BCM46_D_128A
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM46_E
  `define DW_AXI_A2X_RM_BCM46_E `i_axi_a2x_2_DW_AXI_A2X_RM_BCM46_E
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM46_F
  `define DW_AXI_A2X_RM_BCM46_F `i_axi_a2x_2_DW_AXI_A2X_RM_BCM46_F
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM46_X
  `define DW_AXI_A2X_RM_BCM46_X `i_axi_a2x_2_DW_AXI_A2X_RM_BCM46_X
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM47
  `define DW_AXI_A2X_RM_BCM47 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM47
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM48
  `define DW_AXI_A2X_RM_BCM48 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM48
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM48_DM
  `define DW_AXI_A2X_RM_BCM48_DM `i_axi_a2x_2_DW_AXI_A2X_RM_BCM48_DM
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM48_SV
  `define DW_AXI_A2X_RM_BCM48_SV `i_axi_a2x_2_DW_AXI_A2X_RM_BCM48_SV
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM49
  `define DW_AXI_A2X_RM_BCM49 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM49
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM49_SV
  `define DW_AXI_A2X_RM_BCM49_SV `i_axi_a2x_2_DW_AXI_A2X_RM_BCM49_SV
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM50
  `define DW_AXI_A2X_RM_BCM50 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM50
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM51
  `define DW_AXI_A2X_RM_BCM51 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM51
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM52
  `define DW_AXI_A2X_RM_BCM52 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM52
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM53
  `define DW_AXI_A2X_RM_BCM53 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM53
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM54
  `define DW_AXI_A2X_RM_BCM54 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM54
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM55
  `define DW_AXI_A2X_RM_BCM55 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM55
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM55_C
  `define DW_AXI_A2X_RM_BCM55_C `i_axi_a2x_2_DW_AXI_A2X_RM_BCM55_C
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM56
  `define DW_AXI_A2X_RM_BCM56 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM56
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM57
  `define DW_AXI_A2X_RM_BCM57 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM57
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM57_ATV
  `define DW_AXI_A2X_RM_BCM57_ATV `i_axi_a2x_2_DW_AXI_A2X_RM_BCM57_ATV
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM58
  `define DW_AXI_A2X_RM_BCM58 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM58
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM58_ATV
  `define DW_AXI_A2X_RM_BCM58_ATV `i_axi_a2x_2_DW_AXI_A2X_RM_BCM58_ATV
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM59
  `define DW_AXI_A2X_RM_BCM59 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM59
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM60
  `define DW_AXI_A2X_RM_BCM60 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM60
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM62
  `define DW_AXI_A2X_RM_BCM62 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM62
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM63
  `define DW_AXI_A2X_RM_BCM63 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM63
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM64
  `define DW_AXI_A2X_RM_BCM64 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM64
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM64_TD
  `define DW_AXI_A2X_RM_BCM64_TD `i_axi_a2x_2_DW_AXI_A2X_RM_BCM64_TD
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM65
  `define DW_AXI_A2X_RM_BCM65 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM65
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM65_ATV
  `define DW_AXI_A2X_RM_BCM65_ATV `i_axi_a2x_2_DW_AXI_A2X_RM_BCM65_ATV
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM65_TD
  `define DW_AXI_A2X_RM_BCM65_TD `i_axi_a2x_2_DW_AXI_A2X_RM_BCM65_TD
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM66
  `define DW_AXI_A2X_RM_BCM66 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM66
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM66_ATV
  `define DW_AXI_A2X_RM_BCM66_ATV `i_axi_a2x_2_DW_AXI_A2X_RM_BCM66_ATV
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM66_DMS
  `define DW_AXI_A2X_RM_BCM66_DMS `i_axi_a2x_2_DW_AXI_A2X_RM_BCM66_DMS
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM66_DMS_ATV
  `define DW_AXI_A2X_RM_BCM66_DMS_ATV `i_axi_a2x_2_DW_AXI_A2X_RM_BCM66_DMS_ATV
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM66_EFES
  `define DW_AXI_A2X_RM_BCM66_EFES `i_axi_a2x_2_DW_AXI_A2X_RM_BCM66_EFES
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM66_PR
  `define DW_AXI_A2X_RM_BCM66_PR `i_axi_a2x_2_DW_AXI_A2X_RM_BCM66_PR
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM66_WAE
  `define DW_AXI_A2X_RM_BCM66_WAE `i_axi_a2x_2_DW_AXI_A2X_RM_BCM66_WAE
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM66_WAE_ATV
  `define DW_AXI_A2X_RM_BCM66_WAE_ATV `i_axi_a2x_2_DW_AXI_A2X_RM_BCM66_WAE_ATV
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM68_63_7_0
  `define DW_AXI_A2X_RM_BCM68_63_7_0 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM68_63_7_0
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM69_63_7_0
  `define DW_AXI_A2X_RM_BCM69_63_7_0 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM69_63_7_0
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM70_63_7_0_0
  `define DW_AXI_A2X_RM_BCM70_63_7_0_0 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM70_63_7_0_0
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM71
  `define DW_AXI_A2X_RM_BCM71 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM71
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM72
  `define DW_AXI_A2X_RM_BCM72 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM72
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM74
  `define DW_AXI_A2X_RM_BCM74 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM74
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM76
  `define DW_AXI_A2X_RM_BCM76 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM76
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM77
  `define DW_AXI_A2X_RM_BCM77 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM77
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM78
  `define DW_AXI_A2X_RM_BCM78 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM78
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM79
  `define DW_AXI_A2X_RM_BCM79 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM79
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM79_MO
  `define DW_AXI_A2X_RM_BCM79_MO `i_axi_a2x_2_DW_AXI_A2X_RM_BCM79_MO
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM83_GEN
  `define DW_AXI_A2X_RM_BCM83_GEN `i_axi_a2x_2_DW_AXI_A2X_RM_BCM83_GEN
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM84_MON
  `define DW_AXI_A2X_RM_BCM84_MON `i_axi_a2x_2_DW_AXI_A2X_RM_BCM84_MON
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM85
  `define DW_AXI_A2X_RM_BCM85 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM85
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM86
  `define DW_AXI_A2X_RM_BCM86 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM86
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM87
  `define DW_AXI_A2X_RM_BCM87 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM87
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM90
  `define DW_AXI_A2X_RM_BCM90 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM90
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM91
  `define DW_AXI_A2X_RM_BCM91 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM91
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM92
  `define DW_AXI_A2X_RM_BCM92 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM92
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM92_AD
  `define DW_AXI_A2X_RM_BCM92_AD `i_axi_a2x_2_DW_AXI_A2X_RM_BCM92_AD
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM92_AD_DO
  `define DW_AXI_A2X_RM_BCM92_AD_DO `i_axi_a2x_2_DW_AXI_A2X_RM_BCM92_AD_DO
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM92_RD
  `define DW_AXI_A2X_RM_BCM92_RD `i_axi_a2x_2_DW_AXI_A2X_RM_BCM92_RD
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM92_RD_AD
  `define DW_AXI_A2X_RM_BCM92_RD_AD `i_axi_a2x_2_DW_AXI_A2X_RM_BCM92_RD_AD
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM92_RD_AD_DO
  `define DW_AXI_A2X_RM_BCM92_RD_AD_DO `i_axi_a2x_2_DW_AXI_A2X_RM_BCM92_RD_AD_DO
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM92_RD_DO
  `define DW_AXI_A2X_RM_BCM92_RD_DO `i_axi_a2x_2_DW_AXI_A2X_RM_BCM92_RD_DO
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM93
  `define DW_AXI_A2X_RM_BCM93 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM93
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM93_NDSVA
  `define DW_AXI_A2X_RM_BCM93_NDSVA `i_axi_a2x_2_DW_AXI_A2X_RM_BCM93_NDSVA
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM94
  `define DW_AXI_A2X_RM_BCM94 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM94
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM95
  `define DW_AXI_A2X_RM_BCM95 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM95
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM95_E
  `define DW_AXI_A2X_RM_BCM95_E `i_axi_a2x_2_DW_AXI_A2X_RM_BCM95_E
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM95_I
  `define DW_AXI_A2X_RM_BCM95_I `i_axi_a2x_2_DW_AXI_A2X_RM_BCM95_I
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM95_IE
  `define DW_AXI_A2X_RM_BCM95_IE `i_axi_a2x_2_DW_AXI_A2X_RM_BCM95_IE
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM95_NE
  `define DW_AXI_A2X_RM_BCM95_NE `i_axi_a2x_2_DW_AXI_A2X_RM_BCM95_NE
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM95_NE_E
  `define DW_AXI_A2X_RM_BCM95_NE_E `i_axi_a2x_2_DW_AXI_A2X_RM_BCM95_NE_E
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM95_NE_I
  `define DW_AXI_A2X_RM_BCM95_NE_I `i_axi_a2x_2_DW_AXI_A2X_RM_BCM95_NE_I
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM95_NE_IE
  `define DW_AXI_A2X_RM_BCM95_NE_IE `i_axi_a2x_2_DW_AXI_A2X_RM_BCM95_NE_IE
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM98
  `define DW_AXI_A2X_RM_BCM98 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM98
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM99
  `define DW_AXI_A2X_RM_BCM99 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM99
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM99_3
  `define DW_AXI_A2X_RM_BCM99_3 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM99_3
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM99_4
  `define DW_AXI_A2X_RM_BCM99_4 `i_axi_a2x_2_DW_AXI_A2X_RM_BCM99_4
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BCM99_N
  `define DW_AXI_A2X_RM_BCM99_N `i_axi_a2x_2_DW_AXI_A2X_RM_BCM99_N
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BVM01
  `define DW_AXI_A2X_RM_BVM01 `i_axi_a2x_2_DW_AXI_A2X_RM_BVM01
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_BVM02
  `define DW_AXI_A2X_RM_BVM02 `i_axi_a2x_2_DW_AXI_A2X_RM_BVM02
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_SVA01
  `define DW_AXI_A2X_RM_SVA01 `i_axi_a2x_2_DW_AXI_A2X_RM_SVA01
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_SVA02
  `define DW_AXI_A2X_RM_SVA02 `i_axi_a2x_2_DW_AXI_A2X_RM_SVA02
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_SVA03
  `define DW_AXI_A2X_RM_SVA03 `i_axi_a2x_2_DW_AXI_A2X_RM_SVA03
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_SVA04
  `define DW_AXI_A2X_RM_SVA04 `i_axi_a2x_2_DW_AXI_A2X_RM_SVA04
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_SVA05
  `define DW_AXI_A2X_RM_SVA05 `i_axi_a2x_2_DW_AXI_A2X_RM_SVA05
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_SVA06
  `define DW_AXI_A2X_RM_SVA06 `i_axi_a2x_2_DW_AXI_A2X_RM_SVA06
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_SVA07
  `define DW_AXI_A2X_RM_SVA07 `i_axi_a2x_2_DW_AXI_A2X_RM_SVA07
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_SVA08
  `define DW_AXI_A2X_RM_SVA08 `i_axi_a2x_2_DW_AXI_A2X_RM_SVA08
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_SVA09
  `define DW_AXI_A2X_RM_SVA09 `i_axi_a2x_2_DW_AXI_A2X_RM_SVA09
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_SVA10
  `define DW_AXI_A2X_RM_SVA10 `i_axi_a2x_2_DW_AXI_A2X_RM_SVA10
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_SVA11
  `define DW_AXI_A2X_RM_SVA11 `i_axi_a2x_2_DW_AXI_A2X_RM_SVA11
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_SVA12_A
  `define DW_AXI_A2X_RM_SVA12_A `i_axi_a2x_2_DW_AXI_A2X_RM_SVA12_A
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_SVA12_B
  `define DW_AXI_A2X_RM_SVA12_B `i_axi_a2x_2_DW_AXI_A2X_RM_SVA12_B
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_SVA12_C
  `define DW_AXI_A2X_RM_SVA12_C `i_axi_a2x_2_DW_AXI_A2X_RM_SVA12_C
`endif 

`ifdef i_axi_a2x_2_DW_AXI_A2X_RM_SVA99
  `define DW_AXI_A2X_RM_SVA99 `i_axi_a2x_2_DW_AXI_A2X_RM_SVA99
`endif 

`ifdef i_axi_a2x_2___GUARD__DW_AXI_A2X_ALL_INCLUDES__VH__
  `define __GUARD__DW_AXI_A2X_ALL_INCLUDES__VH__ `i_axi_a2x_2___GUARD__DW_AXI_A2X_ALL_INCLUDES__VH__
`endif 

`ifdef i_axi_a2x_2_cb_dummy_parameter_definition
  `define cb_dummy_parameter_definition `i_axi_a2x_2_cb_dummy_parameter_definition
`endif 

