//##########################################################
// Generated undef unprefix file for workspace: DW_axi
//##########################################################

`ifdef __GUARD__DW_AXI_CC_CONSTANTS__VH__
  `undef __GUARD__DW_AXI_CC_CONSTANTS__VH__
`endif 

`ifdef AXI_USE_RANDOM_SEED
  `undef AXI_USE_RANDOM_SEED
`endif 

`ifdef AXI_SEED
  `undef AXI_SEED
`endif 

`ifdef USE_FOUNDATION
  `undef USE_FOUNDATION
`endif 

`ifdef AXI_DW
  `undef AXI_DW
`endif 

`ifdef AXI_AW
  `undef AXI_AW
`endif 

`ifdef AXI_AW_64
  `undef AXI_AW_64
`endif 

`ifdef AXI_NUM_MASTERS
  `undef AXI_NUM_MASTERS
`endif 

`ifdef AXI_NUM_MASTERS_1
  `undef AXI_NUM_MASTERS_1
`endif 

`ifdef AXI_HAS_BICMD
  `undef AXI_HAS_BICMD
`endif 

`ifdef AXI_EN_MULTI_TILE_DLOCK_AVOID
  `undef AXI_EN_MULTI_TILE_DLOCK_AVOID
`endif 

`ifdef AXI_NUM_SYS_MASTERS
  `undef AXI_NUM_SYS_MASTERS
`endif 

`ifdef AXI_NUM_SLAVES
  `undef AXI_NUM_SLAVES
`endif 

`ifdef AXI_LOG2_NS
  `undef AXI_LOG2_NS
`endif 

`ifdef AXI_LOG2_NM
  `undef AXI_LOG2_NM
`endif 

`ifdef AXI_LOG2_LCL_NMP1
  `undef AXI_LOG2_LCL_NMP1
`endif 

`ifdef AXI_LOG2_LCL_NM
  `undef AXI_LOG2_LCL_NM
`endif 

`ifdef AXI_LOG2_NSP1
  `undef AXI_LOG2_NSP1
`endif 

`ifdef AXI_NSP1
  `undef AXI_NSP1
`endif 

`ifdef AXI_LOG2_NSP2
  `undef AXI_LOG2_NSP2
`endif 

`ifdef AXI_MIDW
  `undef AXI_MIDW
`endif 

`ifdef AXI_POW2_MIDW
  `undef AXI_POW2_MIDW
`endif 

`ifdef AXI_SIDW
  `undef AXI_SIDW
`endif 

`ifdef AXI_BLW
  `undef AXI_BLW
`endif 

`ifdef AXI_HAS_TZ_SUPPORT
  `undef AXI_HAS_TZ_SUPPORT
`endif 

`ifdef AXI_TZ_SUPPORT
  `undef AXI_TZ_SUPPORT
`endif 

`ifdef AXI_REMAP_EN
  `undef AXI_REMAP_EN
`endif 

`ifdef AXI_REMAP
  `undef AXI_REMAP
`endif 

`ifdef AXI_HAS_XDCDR
  `undef AXI_HAS_XDCDR
`endif 

`ifdef AXI_XDCDR
  `undef AXI_XDCDR
`endif 

`ifdef AXI_TEST_XDCDR
  `undef AXI_TEST_XDCDR
`endif 

`ifdef AXI_INITIAL_LOCKDOWN
  `undef AXI_INITIAL_LOCKDOWN
`endif 

`ifdef AXI_HAS_LOCKING
  `undef AXI_HAS_LOCKING
`endif 

`ifdef AXI_LOCKING
  `undef AXI_LOCKING
`endif 

`ifdef AXI_LOWPWR_HS_IF
  `undef AXI_LOWPWR_HS_IF
`endif 

`ifdef AXI_LOWPWR_NOPX_CNT
  `undef AXI_LOWPWR_NOPX_CNT
`endif 

`ifdef AXI_LOG2_LOWPWR_NOPX_CNT
  `undef AXI_LOG2_LOWPWR_NOPX_CNT
`endif 

`ifdef AXI_INTERFACE_TYPE
  `undef AXI_INTERFACE_TYPE
`endif 

`ifdef AXI_HAS_AXI4
  `undef AXI_HAS_AXI4
`endif 

`ifdef AXI_HAS_QOS
  `undef AXI_HAS_QOS
`endif 

`ifdef AXI_DLOCK_NOTIFY_EN
  `undef AXI_DLOCK_NOTIFY_EN
`endif 

`ifdef AXI_DLOCK_TIMEOUT
  `undef AXI_DLOCK_TIMEOUT
`endif 

`ifdef AXI_LOG2_DLOCK_TIMEOUT_P1
  `undef AXI_LOG2_DLOCK_TIMEOUT_P1
`endif 

`ifdef AXI_AR_TMO
  `undef AXI_AR_TMO
`endif 

`ifdef AXI_AW_TMO
  `undef AXI_AW_TMO
`endif 

`ifdef AXI_W_TMO
  `undef AXI_W_TMO
`endif 

`ifdef AXI_R_TMO
  `undef AXI_R_TMO
`endif 

`ifdef AXI_B_TMO
  `undef AXI_B_TMO
`endif 

`ifdef AXI_AR_PL_ARB
  `undef AXI_AR_PL_ARB
`endif 

`ifdef AXI_AW_PL_ARB
  `undef AXI_AW_PL_ARB
`endif 

`ifdef AXI_R_PL_ARB
  `undef AXI_R_PL_ARB
`endif 

`ifdef AXI_W_PL_ARB
  `undef AXI_W_PL_ARB
`endif 

`ifdef AXI_B_PL_ARB
  `undef AXI_B_PL_ARB
`endif 

`ifdef AXI_ENCRYPT
  `undef AXI_ENCRYPT
`endif 

`ifdef AXI_MST_PRIORITY_W
  `undef AXI_MST_PRIORITY_W
`endif 

`ifdef AXI_SLV_PRIORITY_W
  `undef AXI_SLV_PRIORITY_W
`endif 

`ifdef AXI_REG_AW_W_PATHS
  `undef AXI_REG_AW_W_PATHS
`endif 

`ifdef AXI_MAX_UIDA
  `undef AXI_MAX_UIDA
`endif 

`ifdef AXI_HAS_LEGAL_ADDR_OVRLP_VAL
  `undef AXI_HAS_LEGAL_ADDR_OVRLP_VAL
`endif 

`ifdef AXI_HAS_LEGAL_ADDR_OVRLP
  `undef AXI_HAS_LEGAL_ADDR_OVRLP
`endif 

`ifdef AXI_VLD_RDY_PARITY_PROT
  `undef AXI_VLD_RDY_PARITY_PROT
`endif 

`ifdef AXI_VLD_RDY_PARITY_MODE
  `undef AXI_VLD_RDY_PARITY_MODE
`endif 

`ifdef AXI_HAS_EVEN_PARITY
  `undef AXI_HAS_EVEN_PARITY
`endif 

`ifdef IFX_RULE_SETUP
  `undef IFX_RULE_SETUP
`endif 

`ifdef AXI_INTF_PAR_EN
  `undef AXI_INTF_PAR_EN
`endif 

`ifdef AXI_INTF_PARITY_MODE
  `undef AXI_INTF_PARITY_MODE
`endif 

`ifdef AXI_MAX_SBW
  `undef AXI_MAX_SBW
`endif 

`ifdef AXI_HAS_AWSB
  `undef AXI_HAS_AWSB
`endif 

`ifdef AXI_INC_AWSB
  `undef AXI_INC_AWSB
`endif 

`ifdef AXI_AW_SBW
  `undef AXI_AW_SBW
`endif 

`ifdef AXI_HAS_WSB
  `undef AXI_HAS_WSB
`endif 

`ifdef AXI_INC_WSB
  `undef AXI_INC_WSB
`endif 

`ifdef AXI_W_SBW
  `undef AXI_W_SBW
`endif 

`ifdef AXI_HAS_BSB
  `undef AXI_HAS_BSB
`endif 

`ifdef AXI_INC_BSB
  `undef AXI_INC_BSB
`endif 

`ifdef AXI_B_SBW
  `undef AXI_B_SBW
`endif 

`ifdef AXI_HAS_ARSB
  `undef AXI_HAS_ARSB
`endif 

`ifdef AXI_INC_ARSB
  `undef AXI_INC_ARSB
`endif 

`ifdef AXI_AR_SBW
  `undef AXI_AR_SBW
`endif 

`ifdef AXI_HAS_RSB
  `undef AXI_HAS_RSB
`endif 

`ifdef AXI_INC_RSB
  `undef AXI_INC_RSB
`endif 

`ifdef AXI_R_SBW
  `undef AXI_R_SBW
`endif 

`ifdef AXI_NV_S0_BY_M1
  `undef AXI_NV_S0_BY_M1
`endif 

`ifdef AXI_NV_S0_BY_M2
  `undef AXI_NV_S0_BY_M2
`endif 

`ifdef AXI_NV_S0_BY_M3
  `undef AXI_NV_S0_BY_M3
`endif 

`ifdef AXI_NV_S0_BY_M4
  `undef AXI_NV_S0_BY_M4
`endif 

`ifdef AXI_NV_S0_BY_M5
  `undef AXI_NV_S0_BY_M5
`endif 

`ifdef AXI_NV_S0_BY_M6
  `undef AXI_NV_S0_BY_M6
`endif 

`ifdef AXI_NV_S0_BY_M7
  `undef AXI_NV_S0_BY_M7
`endif 

`ifdef AXI_NV_S0_BY_M8
  `undef AXI_NV_S0_BY_M8
`endif 

`ifdef AXI_NV_S0_BY_M9
  `undef AXI_NV_S0_BY_M9
`endif 

`ifdef AXI_NV_S0_BY_M10
  `undef AXI_NV_S0_BY_M10
`endif 

`ifdef AXI_NV_S0_BY_M11
  `undef AXI_NV_S0_BY_M11
`endif 

`ifdef AXI_NV_S0_BY_M12
  `undef AXI_NV_S0_BY_M12
`endif 

`ifdef AXI_NV_S0_BY_M13
  `undef AXI_NV_S0_BY_M13
`endif 

`ifdef AXI_NV_S0_BY_M14
  `undef AXI_NV_S0_BY_M14
`endif 

`ifdef AXI_NV_S0_BY_M15
  `undef AXI_NV_S0_BY_M15
`endif 

`ifdef AXI_NV_S0_BY_M16
  `undef AXI_NV_S0_BY_M16
`endif 

`ifdef AXI_NV_S1_BY_M1
  `undef AXI_NV_S1_BY_M1
`endif 

`ifdef AXI_NV_S1_BY_M2
  `undef AXI_NV_S1_BY_M2
`endif 

`ifdef AXI_NV_S1_BY_M3
  `undef AXI_NV_S1_BY_M3
`endif 

`ifdef AXI_NV_S1_BY_M4
  `undef AXI_NV_S1_BY_M4
`endif 

`ifdef AXI_NV_S1_BY_M5
  `undef AXI_NV_S1_BY_M5
`endif 

`ifdef AXI_NV_S1_BY_M6
  `undef AXI_NV_S1_BY_M6
`endif 

`ifdef AXI_NV_S1_BY_M7
  `undef AXI_NV_S1_BY_M7
`endif 

`ifdef AXI_NV_S1_BY_M8
  `undef AXI_NV_S1_BY_M8
`endif 

`ifdef AXI_NV_S1_BY_M9
  `undef AXI_NV_S1_BY_M9
`endif 

`ifdef AXI_NV_S1_BY_M10
  `undef AXI_NV_S1_BY_M10
`endif 

`ifdef AXI_NV_S1_BY_M11
  `undef AXI_NV_S1_BY_M11
`endif 

`ifdef AXI_NV_S1_BY_M12
  `undef AXI_NV_S1_BY_M12
`endif 

`ifdef AXI_NV_S1_BY_M13
  `undef AXI_NV_S1_BY_M13
`endif 

`ifdef AXI_NV_S1_BY_M14
  `undef AXI_NV_S1_BY_M14
`endif 

`ifdef AXI_NV_S1_BY_M15
  `undef AXI_NV_S1_BY_M15
`endif 

`ifdef AXI_NV_S1_BY_M16
  `undef AXI_NV_S1_BY_M16
`endif 

`ifdef AXI_NV_S2_BY_M1
  `undef AXI_NV_S2_BY_M1
`endif 

`ifdef AXI_NV_S2_BY_M2
  `undef AXI_NV_S2_BY_M2
`endif 

`ifdef AXI_NV_S2_BY_M3
  `undef AXI_NV_S2_BY_M3
`endif 

`ifdef AXI_NV_S2_BY_M4
  `undef AXI_NV_S2_BY_M4
`endif 

`ifdef AXI_NV_S2_BY_M5
  `undef AXI_NV_S2_BY_M5
`endif 

`ifdef AXI_NV_S2_BY_M6
  `undef AXI_NV_S2_BY_M6
`endif 

`ifdef AXI_NV_S2_BY_M7
  `undef AXI_NV_S2_BY_M7
`endif 

`ifdef AXI_NV_S2_BY_M8
  `undef AXI_NV_S2_BY_M8
`endif 

`ifdef AXI_NV_S2_BY_M9
  `undef AXI_NV_S2_BY_M9
`endif 

`ifdef AXI_NV_S2_BY_M10
  `undef AXI_NV_S2_BY_M10
`endif 

`ifdef AXI_NV_S2_BY_M11
  `undef AXI_NV_S2_BY_M11
`endif 

`ifdef AXI_NV_S2_BY_M12
  `undef AXI_NV_S2_BY_M12
`endif 

`ifdef AXI_NV_S2_BY_M13
  `undef AXI_NV_S2_BY_M13
`endif 

`ifdef AXI_NV_S2_BY_M14
  `undef AXI_NV_S2_BY_M14
`endif 

`ifdef AXI_NV_S2_BY_M15
  `undef AXI_NV_S2_BY_M15
`endif 

`ifdef AXI_NV_S2_BY_M16
  `undef AXI_NV_S2_BY_M16
`endif 

`ifdef AXI_NV_S3_BY_M1
  `undef AXI_NV_S3_BY_M1
`endif 

`ifdef AXI_NV_S3_BY_M2
  `undef AXI_NV_S3_BY_M2
`endif 

`ifdef AXI_NV_S3_BY_M3
  `undef AXI_NV_S3_BY_M3
`endif 

`ifdef AXI_NV_S3_BY_M4
  `undef AXI_NV_S3_BY_M4
`endif 

`ifdef AXI_NV_S3_BY_M5
  `undef AXI_NV_S3_BY_M5
`endif 

`ifdef AXI_NV_S3_BY_M6
  `undef AXI_NV_S3_BY_M6
`endif 

`ifdef AXI_NV_S3_BY_M7
  `undef AXI_NV_S3_BY_M7
`endif 

`ifdef AXI_NV_S3_BY_M8
  `undef AXI_NV_S3_BY_M8
`endif 

`ifdef AXI_NV_S3_BY_M9
  `undef AXI_NV_S3_BY_M9
`endif 

`ifdef AXI_NV_S3_BY_M10
  `undef AXI_NV_S3_BY_M10
`endif 

`ifdef AXI_NV_S3_BY_M11
  `undef AXI_NV_S3_BY_M11
`endif 

`ifdef AXI_NV_S3_BY_M12
  `undef AXI_NV_S3_BY_M12
`endif 

`ifdef AXI_NV_S3_BY_M13
  `undef AXI_NV_S3_BY_M13
`endif 

`ifdef AXI_NV_S3_BY_M14
  `undef AXI_NV_S3_BY_M14
`endif 

`ifdef AXI_NV_S3_BY_M15
  `undef AXI_NV_S3_BY_M15
`endif 

`ifdef AXI_NV_S3_BY_M16
  `undef AXI_NV_S3_BY_M16
`endif 

`ifdef AXI_NV_S4_BY_M1
  `undef AXI_NV_S4_BY_M1
`endif 

`ifdef AXI_NV_S4_BY_M2
  `undef AXI_NV_S4_BY_M2
`endif 

`ifdef AXI_NV_S4_BY_M3
  `undef AXI_NV_S4_BY_M3
`endif 

`ifdef AXI_NV_S4_BY_M4
  `undef AXI_NV_S4_BY_M4
`endif 

`ifdef AXI_NV_S4_BY_M5
  `undef AXI_NV_S4_BY_M5
`endif 

`ifdef AXI_NV_S4_BY_M6
  `undef AXI_NV_S4_BY_M6
`endif 

`ifdef AXI_NV_S4_BY_M7
  `undef AXI_NV_S4_BY_M7
`endif 

`ifdef AXI_NV_S4_BY_M8
  `undef AXI_NV_S4_BY_M8
`endif 

`ifdef AXI_NV_S4_BY_M9
  `undef AXI_NV_S4_BY_M9
`endif 

`ifdef AXI_NV_S4_BY_M10
  `undef AXI_NV_S4_BY_M10
`endif 

`ifdef AXI_NV_S4_BY_M11
  `undef AXI_NV_S4_BY_M11
`endif 

`ifdef AXI_NV_S4_BY_M12
  `undef AXI_NV_S4_BY_M12
`endif 

`ifdef AXI_NV_S4_BY_M13
  `undef AXI_NV_S4_BY_M13
`endif 

`ifdef AXI_NV_S4_BY_M14
  `undef AXI_NV_S4_BY_M14
`endif 

`ifdef AXI_NV_S4_BY_M15
  `undef AXI_NV_S4_BY_M15
`endif 

`ifdef AXI_NV_S4_BY_M16
  `undef AXI_NV_S4_BY_M16
`endif 

`ifdef AXI_NV_S5_BY_M1
  `undef AXI_NV_S5_BY_M1
`endif 

`ifdef AXI_NV_S5_BY_M2
  `undef AXI_NV_S5_BY_M2
`endif 

`ifdef AXI_NV_S5_BY_M3
  `undef AXI_NV_S5_BY_M3
`endif 

`ifdef AXI_NV_S5_BY_M4
  `undef AXI_NV_S5_BY_M4
`endif 

`ifdef AXI_NV_S5_BY_M5
  `undef AXI_NV_S5_BY_M5
`endif 

`ifdef AXI_NV_S5_BY_M6
  `undef AXI_NV_S5_BY_M6
`endif 

`ifdef AXI_NV_S5_BY_M7
  `undef AXI_NV_S5_BY_M7
`endif 

`ifdef AXI_NV_S5_BY_M8
  `undef AXI_NV_S5_BY_M8
`endif 

`ifdef AXI_NV_S5_BY_M9
  `undef AXI_NV_S5_BY_M9
`endif 

`ifdef AXI_NV_S5_BY_M10
  `undef AXI_NV_S5_BY_M10
`endif 

`ifdef AXI_NV_S5_BY_M11
  `undef AXI_NV_S5_BY_M11
`endif 

`ifdef AXI_NV_S5_BY_M12
  `undef AXI_NV_S5_BY_M12
`endif 

`ifdef AXI_NV_S5_BY_M13
  `undef AXI_NV_S5_BY_M13
`endif 

`ifdef AXI_NV_S5_BY_M14
  `undef AXI_NV_S5_BY_M14
`endif 

`ifdef AXI_NV_S5_BY_M15
  `undef AXI_NV_S5_BY_M15
`endif 

`ifdef AXI_NV_S5_BY_M16
  `undef AXI_NV_S5_BY_M16
`endif 

`ifdef AXI_NV_S6_BY_M1
  `undef AXI_NV_S6_BY_M1
`endif 

`ifdef AXI_NV_S6_BY_M2
  `undef AXI_NV_S6_BY_M2
`endif 

`ifdef AXI_NV_S6_BY_M3
  `undef AXI_NV_S6_BY_M3
`endif 

`ifdef AXI_NV_S6_BY_M4
  `undef AXI_NV_S6_BY_M4
`endif 

`ifdef AXI_NV_S6_BY_M5
  `undef AXI_NV_S6_BY_M5
`endif 

`ifdef AXI_NV_S6_BY_M6
  `undef AXI_NV_S6_BY_M6
`endif 

`ifdef AXI_NV_S6_BY_M7
  `undef AXI_NV_S6_BY_M7
`endif 

`ifdef AXI_NV_S6_BY_M8
  `undef AXI_NV_S6_BY_M8
`endif 

`ifdef AXI_NV_S6_BY_M9
  `undef AXI_NV_S6_BY_M9
`endif 

`ifdef AXI_NV_S6_BY_M10
  `undef AXI_NV_S6_BY_M10
`endif 

`ifdef AXI_NV_S6_BY_M11
  `undef AXI_NV_S6_BY_M11
`endif 

`ifdef AXI_NV_S6_BY_M12
  `undef AXI_NV_S6_BY_M12
`endif 

`ifdef AXI_NV_S6_BY_M13
  `undef AXI_NV_S6_BY_M13
`endif 

`ifdef AXI_NV_S6_BY_M14
  `undef AXI_NV_S6_BY_M14
`endif 

`ifdef AXI_NV_S6_BY_M15
  `undef AXI_NV_S6_BY_M15
`endif 

`ifdef AXI_NV_S6_BY_M16
  `undef AXI_NV_S6_BY_M16
`endif 

`ifdef AXI_NV_S7_BY_M1
  `undef AXI_NV_S7_BY_M1
`endif 

`ifdef AXI_NV_S7_BY_M2
  `undef AXI_NV_S7_BY_M2
`endif 

`ifdef AXI_NV_S7_BY_M3
  `undef AXI_NV_S7_BY_M3
`endif 

`ifdef AXI_NV_S7_BY_M4
  `undef AXI_NV_S7_BY_M4
`endif 

`ifdef AXI_NV_S7_BY_M5
  `undef AXI_NV_S7_BY_M5
`endif 

`ifdef AXI_NV_S7_BY_M6
  `undef AXI_NV_S7_BY_M6
`endif 

`ifdef AXI_NV_S7_BY_M7
  `undef AXI_NV_S7_BY_M7
`endif 

`ifdef AXI_NV_S7_BY_M8
  `undef AXI_NV_S7_BY_M8
`endif 

`ifdef AXI_NV_S7_BY_M9
  `undef AXI_NV_S7_BY_M9
`endif 

`ifdef AXI_NV_S7_BY_M10
  `undef AXI_NV_S7_BY_M10
`endif 

`ifdef AXI_NV_S7_BY_M11
  `undef AXI_NV_S7_BY_M11
`endif 

`ifdef AXI_NV_S7_BY_M12
  `undef AXI_NV_S7_BY_M12
`endif 

`ifdef AXI_NV_S7_BY_M13
  `undef AXI_NV_S7_BY_M13
`endif 

`ifdef AXI_NV_S7_BY_M14
  `undef AXI_NV_S7_BY_M14
`endif 

`ifdef AXI_NV_S7_BY_M15
  `undef AXI_NV_S7_BY_M15
`endif 

`ifdef AXI_NV_S7_BY_M16
  `undef AXI_NV_S7_BY_M16
`endif 

`ifdef AXI_NV_S8_BY_M1
  `undef AXI_NV_S8_BY_M1
`endif 

`ifdef AXI_NV_S8_BY_M2
  `undef AXI_NV_S8_BY_M2
`endif 

`ifdef AXI_NV_S8_BY_M3
  `undef AXI_NV_S8_BY_M3
`endif 

`ifdef AXI_NV_S8_BY_M4
  `undef AXI_NV_S8_BY_M4
`endif 

`ifdef AXI_NV_S8_BY_M5
  `undef AXI_NV_S8_BY_M5
`endif 

`ifdef AXI_NV_S8_BY_M6
  `undef AXI_NV_S8_BY_M6
`endif 

`ifdef AXI_NV_S8_BY_M7
  `undef AXI_NV_S8_BY_M7
`endif 

`ifdef AXI_NV_S8_BY_M8
  `undef AXI_NV_S8_BY_M8
`endif 

`ifdef AXI_NV_S8_BY_M9
  `undef AXI_NV_S8_BY_M9
`endif 

`ifdef AXI_NV_S8_BY_M10
  `undef AXI_NV_S8_BY_M10
`endif 

`ifdef AXI_NV_S8_BY_M11
  `undef AXI_NV_S8_BY_M11
`endif 

`ifdef AXI_NV_S8_BY_M12
  `undef AXI_NV_S8_BY_M12
`endif 

`ifdef AXI_NV_S8_BY_M13
  `undef AXI_NV_S8_BY_M13
`endif 

`ifdef AXI_NV_S8_BY_M14
  `undef AXI_NV_S8_BY_M14
`endif 

`ifdef AXI_NV_S8_BY_M15
  `undef AXI_NV_S8_BY_M15
`endif 

`ifdef AXI_NV_S8_BY_M16
  `undef AXI_NV_S8_BY_M16
`endif 

`ifdef AXI_NV_S9_BY_M1
  `undef AXI_NV_S9_BY_M1
`endif 

`ifdef AXI_NV_S9_BY_M2
  `undef AXI_NV_S9_BY_M2
`endif 

`ifdef AXI_NV_S9_BY_M3
  `undef AXI_NV_S9_BY_M3
`endif 

`ifdef AXI_NV_S9_BY_M4
  `undef AXI_NV_S9_BY_M4
`endif 

`ifdef AXI_NV_S9_BY_M5
  `undef AXI_NV_S9_BY_M5
`endif 

`ifdef AXI_NV_S9_BY_M6
  `undef AXI_NV_S9_BY_M6
`endif 

`ifdef AXI_NV_S9_BY_M7
  `undef AXI_NV_S9_BY_M7
`endif 

`ifdef AXI_NV_S9_BY_M8
  `undef AXI_NV_S9_BY_M8
`endif 

`ifdef AXI_NV_S9_BY_M9
  `undef AXI_NV_S9_BY_M9
`endif 

`ifdef AXI_NV_S9_BY_M10
  `undef AXI_NV_S9_BY_M10
`endif 

`ifdef AXI_NV_S9_BY_M11
  `undef AXI_NV_S9_BY_M11
`endif 

`ifdef AXI_NV_S9_BY_M12
  `undef AXI_NV_S9_BY_M12
`endif 

`ifdef AXI_NV_S9_BY_M13
  `undef AXI_NV_S9_BY_M13
`endif 

`ifdef AXI_NV_S9_BY_M14
  `undef AXI_NV_S9_BY_M14
`endif 

`ifdef AXI_NV_S9_BY_M15
  `undef AXI_NV_S9_BY_M15
`endif 

`ifdef AXI_NV_S9_BY_M16
  `undef AXI_NV_S9_BY_M16
`endif 

`ifdef AXI_NV_S10_BY_M1
  `undef AXI_NV_S10_BY_M1
`endif 

`ifdef AXI_NV_S10_BY_M2
  `undef AXI_NV_S10_BY_M2
`endif 

`ifdef AXI_NV_S10_BY_M3
  `undef AXI_NV_S10_BY_M3
`endif 

`ifdef AXI_NV_S10_BY_M4
  `undef AXI_NV_S10_BY_M4
`endif 

`ifdef AXI_NV_S10_BY_M5
  `undef AXI_NV_S10_BY_M5
`endif 

`ifdef AXI_NV_S10_BY_M6
  `undef AXI_NV_S10_BY_M6
`endif 

`ifdef AXI_NV_S10_BY_M7
  `undef AXI_NV_S10_BY_M7
`endif 

`ifdef AXI_NV_S10_BY_M8
  `undef AXI_NV_S10_BY_M8
`endif 

`ifdef AXI_NV_S10_BY_M9
  `undef AXI_NV_S10_BY_M9
`endif 

`ifdef AXI_NV_S10_BY_M10
  `undef AXI_NV_S10_BY_M10
`endif 

`ifdef AXI_NV_S10_BY_M11
  `undef AXI_NV_S10_BY_M11
`endif 

`ifdef AXI_NV_S10_BY_M12
  `undef AXI_NV_S10_BY_M12
`endif 

`ifdef AXI_NV_S10_BY_M13
  `undef AXI_NV_S10_BY_M13
`endif 

`ifdef AXI_NV_S10_BY_M14
  `undef AXI_NV_S10_BY_M14
`endif 

`ifdef AXI_NV_S10_BY_M15
  `undef AXI_NV_S10_BY_M15
`endif 

`ifdef AXI_NV_S10_BY_M16
  `undef AXI_NV_S10_BY_M16
`endif 

`ifdef AXI_NV_S11_BY_M1
  `undef AXI_NV_S11_BY_M1
`endif 

`ifdef AXI_NV_S11_BY_M2
  `undef AXI_NV_S11_BY_M2
`endif 

`ifdef AXI_NV_S11_BY_M3
  `undef AXI_NV_S11_BY_M3
`endif 

`ifdef AXI_NV_S11_BY_M4
  `undef AXI_NV_S11_BY_M4
`endif 

`ifdef AXI_NV_S11_BY_M5
  `undef AXI_NV_S11_BY_M5
`endif 

`ifdef AXI_NV_S11_BY_M6
  `undef AXI_NV_S11_BY_M6
`endif 

`ifdef AXI_NV_S11_BY_M7
  `undef AXI_NV_S11_BY_M7
`endif 

`ifdef AXI_NV_S11_BY_M8
  `undef AXI_NV_S11_BY_M8
`endif 

`ifdef AXI_NV_S11_BY_M9
  `undef AXI_NV_S11_BY_M9
`endif 

`ifdef AXI_NV_S11_BY_M10
  `undef AXI_NV_S11_BY_M10
`endif 

`ifdef AXI_NV_S11_BY_M11
  `undef AXI_NV_S11_BY_M11
`endif 

`ifdef AXI_NV_S11_BY_M12
  `undef AXI_NV_S11_BY_M12
`endif 

`ifdef AXI_NV_S11_BY_M13
  `undef AXI_NV_S11_BY_M13
`endif 

`ifdef AXI_NV_S11_BY_M14
  `undef AXI_NV_S11_BY_M14
`endif 

`ifdef AXI_NV_S11_BY_M15
  `undef AXI_NV_S11_BY_M15
`endif 

`ifdef AXI_NV_S11_BY_M16
  `undef AXI_NV_S11_BY_M16
`endif 

`ifdef AXI_NV_S12_BY_M1
  `undef AXI_NV_S12_BY_M1
`endif 

`ifdef AXI_NV_S12_BY_M2
  `undef AXI_NV_S12_BY_M2
`endif 

`ifdef AXI_NV_S12_BY_M3
  `undef AXI_NV_S12_BY_M3
`endif 

`ifdef AXI_NV_S12_BY_M4
  `undef AXI_NV_S12_BY_M4
`endif 

`ifdef AXI_NV_S12_BY_M5
  `undef AXI_NV_S12_BY_M5
`endif 

`ifdef AXI_NV_S12_BY_M6
  `undef AXI_NV_S12_BY_M6
`endif 

`ifdef AXI_NV_S12_BY_M7
  `undef AXI_NV_S12_BY_M7
`endif 

`ifdef AXI_NV_S12_BY_M8
  `undef AXI_NV_S12_BY_M8
`endif 

`ifdef AXI_NV_S12_BY_M9
  `undef AXI_NV_S12_BY_M9
`endif 

`ifdef AXI_NV_S12_BY_M10
  `undef AXI_NV_S12_BY_M10
`endif 

`ifdef AXI_NV_S12_BY_M11
  `undef AXI_NV_S12_BY_M11
`endif 

`ifdef AXI_NV_S12_BY_M12
  `undef AXI_NV_S12_BY_M12
`endif 

`ifdef AXI_NV_S12_BY_M13
  `undef AXI_NV_S12_BY_M13
`endif 

`ifdef AXI_NV_S12_BY_M14
  `undef AXI_NV_S12_BY_M14
`endif 

`ifdef AXI_NV_S12_BY_M15
  `undef AXI_NV_S12_BY_M15
`endif 

`ifdef AXI_NV_S12_BY_M16
  `undef AXI_NV_S12_BY_M16
`endif 

`ifdef AXI_NV_S13_BY_M1
  `undef AXI_NV_S13_BY_M1
`endif 

`ifdef AXI_NV_S13_BY_M2
  `undef AXI_NV_S13_BY_M2
`endif 

`ifdef AXI_NV_S13_BY_M3
  `undef AXI_NV_S13_BY_M3
`endif 

`ifdef AXI_NV_S13_BY_M4
  `undef AXI_NV_S13_BY_M4
`endif 

`ifdef AXI_NV_S13_BY_M5
  `undef AXI_NV_S13_BY_M5
`endif 

`ifdef AXI_NV_S13_BY_M6
  `undef AXI_NV_S13_BY_M6
`endif 

`ifdef AXI_NV_S13_BY_M7
  `undef AXI_NV_S13_BY_M7
`endif 

`ifdef AXI_NV_S13_BY_M8
  `undef AXI_NV_S13_BY_M8
`endif 

`ifdef AXI_NV_S13_BY_M9
  `undef AXI_NV_S13_BY_M9
`endif 

`ifdef AXI_NV_S13_BY_M10
  `undef AXI_NV_S13_BY_M10
`endif 

`ifdef AXI_NV_S13_BY_M11
  `undef AXI_NV_S13_BY_M11
`endif 

`ifdef AXI_NV_S13_BY_M12
  `undef AXI_NV_S13_BY_M12
`endif 

`ifdef AXI_NV_S13_BY_M13
  `undef AXI_NV_S13_BY_M13
`endif 

`ifdef AXI_NV_S13_BY_M14
  `undef AXI_NV_S13_BY_M14
`endif 

`ifdef AXI_NV_S13_BY_M15
  `undef AXI_NV_S13_BY_M15
`endif 

`ifdef AXI_NV_S13_BY_M16
  `undef AXI_NV_S13_BY_M16
`endif 

`ifdef AXI_NV_S14_BY_M1
  `undef AXI_NV_S14_BY_M1
`endif 

`ifdef AXI_NV_S14_BY_M2
  `undef AXI_NV_S14_BY_M2
`endif 

`ifdef AXI_NV_S14_BY_M3
  `undef AXI_NV_S14_BY_M3
`endif 

`ifdef AXI_NV_S14_BY_M4
  `undef AXI_NV_S14_BY_M4
`endif 

`ifdef AXI_NV_S14_BY_M5
  `undef AXI_NV_S14_BY_M5
`endif 

`ifdef AXI_NV_S14_BY_M6
  `undef AXI_NV_S14_BY_M6
`endif 

`ifdef AXI_NV_S14_BY_M7
  `undef AXI_NV_S14_BY_M7
`endif 

`ifdef AXI_NV_S14_BY_M8
  `undef AXI_NV_S14_BY_M8
`endif 

`ifdef AXI_NV_S14_BY_M9
  `undef AXI_NV_S14_BY_M9
`endif 

`ifdef AXI_NV_S14_BY_M10
  `undef AXI_NV_S14_BY_M10
`endif 

`ifdef AXI_NV_S14_BY_M11
  `undef AXI_NV_S14_BY_M11
`endif 

`ifdef AXI_NV_S14_BY_M12
  `undef AXI_NV_S14_BY_M12
`endif 

`ifdef AXI_NV_S14_BY_M13
  `undef AXI_NV_S14_BY_M13
`endif 

`ifdef AXI_NV_S14_BY_M14
  `undef AXI_NV_S14_BY_M14
`endif 

`ifdef AXI_NV_S14_BY_M15
  `undef AXI_NV_S14_BY_M15
`endif 

`ifdef AXI_NV_S14_BY_M16
  `undef AXI_NV_S14_BY_M16
`endif 

`ifdef AXI_NV_S15_BY_M1
  `undef AXI_NV_S15_BY_M1
`endif 

`ifdef AXI_NV_S15_BY_M2
  `undef AXI_NV_S15_BY_M2
`endif 

`ifdef AXI_NV_S15_BY_M3
  `undef AXI_NV_S15_BY_M3
`endif 

`ifdef AXI_NV_S15_BY_M4
  `undef AXI_NV_S15_BY_M4
`endif 

`ifdef AXI_NV_S15_BY_M5
  `undef AXI_NV_S15_BY_M5
`endif 

`ifdef AXI_NV_S15_BY_M6
  `undef AXI_NV_S15_BY_M6
`endif 

`ifdef AXI_NV_S15_BY_M7
  `undef AXI_NV_S15_BY_M7
`endif 

`ifdef AXI_NV_S15_BY_M8
  `undef AXI_NV_S15_BY_M8
`endif 

`ifdef AXI_NV_S15_BY_M9
  `undef AXI_NV_S15_BY_M9
`endif 

`ifdef AXI_NV_S15_BY_M10
  `undef AXI_NV_S15_BY_M10
`endif 

`ifdef AXI_NV_S15_BY_M11
  `undef AXI_NV_S15_BY_M11
`endif 

`ifdef AXI_NV_S15_BY_M12
  `undef AXI_NV_S15_BY_M12
`endif 

`ifdef AXI_NV_S15_BY_M13
  `undef AXI_NV_S15_BY_M13
`endif 

`ifdef AXI_NV_S15_BY_M14
  `undef AXI_NV_S15_BY_M14
`endif 

`ifdef AXI_NV_S15_BY_M15
  `undef AXI_NV_S15_BY_M15
`endif 

`ifdef AXI_NV_S15_BY_M16
  `undef AXI_NV_S15_BY_M16
`endif 

`ifdef AXI_NV_S16_BY_M1
  `undef AXI_NV_S16_BY_M1
`endif 

`ifdef AXI_NV_S16_BY_M2
  `undef AXI_NV_S16_BY_M2
`endif 

`ifdef AXI_NV_S16_BY_M3
  `undef AXI_NV_S16_BY_M3
`endif 

`ifdef AXI_NV_S16_BY_M4
  `undef AXI_NV_S16_BY_M4
`endif 

`ifdef AXI_NV_S16_BY_M5
  `undef AXI_NV_S16_BY_M5
`endif 

`ifdef AXI_NV_S16_BY_M6
  `undef AXI_NV_S16_BY_M6
`endif 

`ifdef AXI_NV_S16_BY_M7
  `undef AXI_NV_S16_BY_M7
`endif 

`ifdef AXI_NV_S16_BY_M8
  `undef AXI_NV_S16_BY_M8
`endif 

`ifdef AXI_NV_S16_BY_M9
  `undef AXI_NV_S16_BY_M9
`endif 

`ifdef AXI_NV_S16_BY_M10
  `undef AXI_NV_S16_BY_M10
`endif 

`ifdef AXI_NV_S16_BY_M11
  `undef AXI_NV_S16_BY_M11
`endif 

`ifdef AXI_NV_S16_BY_M12
  `undef AXI_NV_S16_BY_M12
`endif 

`ifdef AXI_NV_S16_BY_M13
  `undef AXI_NV_S16_BY_M13
`endif 

`ifdef AXI_NV_S16_BY_M14
  `undef AXI_NV_S16_BY_M14
`endif 

`ifdef AXI_NV_S16_BY_M15
  `undef AXI_NV_S16_BY_M15
`endif 

`ifdef AXI_NV_S16_BY_M16
  `undef AXI_NV_S16_BY_M16
`endif 

`ifdef AXI_NV_S1_BY_ANY_M
  `undef AXI_NV_S1_BY_ANY_M
`endif 

`ifdef AXI_NV_S2_BY_ANY_M
  `undef AXI_NV_S2_BY_ANY_M
`endif 

`ifdef AXI_NV_S3_BY_ANY_M
  `undef AXI_NV_S3_BY_ANY_M
`endif 

`ifdef AXI_NV_S4_BY_ANY_M
  `undef AXI_NV_S4_BY_ANY_M
`endif 

`ifdef AXI_NV_S5_BY_ANY_M
  `undef AXI_NV_S5_BY_ANY_M
`endif 

`ifdef AXI_NV_S6_BY_ANY_M
  `undef AXI_NV_S6_BY_ANY_M
`endif 

`ifdef AXI_NV_S7_BY_ANY_M
  `undef AXI_NV_S7_BY_ANY_M
`endif 

`ifdef AXI_NV_S8_BY_ANY_M
  `undef AXI_NV_S8_BY_ANY_M
`endif 

`ifdef AXI_NV_S9_BY_ANY_M
  `undef AXI_NV_S9_BY_ANY_M
`endif 

`ifdef AXI_NV_S10_BY_ANY_M
  `undef AXI_NV_S10_BY_ANY_M
`endif 

`ifdef AXI_NV_S11_BY_ANY_M
  `undef AXI_NV_S11_BY_ANY_M
`endif 

`ifdef AXI_NV_S12_BY_ANY_M
  `undef AXI_NV_S12_BY_ANY_M
`endif 

`ifdef AXI_NV_S13_BY_ANY_M
  `undef AXI_NV_S13_BY_ANY_M
`endif 

`ifdef AXI_NV_S14_BY_ANY_M
  `undef AXI_NV_S14_BY_ANY_M
`endif 

`ifdef AXI_NV_S15_BY_ANY_M
  `undef AXI_NV_S15_BY_ANY_M
`endif 

`ifdef AXI_NV_S16_BY_ANY_M
  `undef AXI_NV_S16_BY_ANY_M
`endif 

`ifdef AXI_BV_S0_BY_M1
  `undef AXI_BV_S0_BY_M1
`endif 

`ifdef AXI_BV_S0_BY_M2
  `undef AXI_BV_S0_BY_M2
`endif 

`ifdef AXI_BV_S0_BY_M3
  `undef AXI_BV_S0_BY_M3
`endif 

`ifdef AXI_BV_S0_BY_M4
  `undef AXI_BV_S0_BY_M4
`endif 

`ifdef AXI_BV_S0_BY_M5
  `undef AXI_BV_S0_BY_M5
`endif 

`ifdef AXI_BV_S0_BY_M6
  `undef AXI_BV_S0_BY_M6
`endif 

`ifdef AXI_BV_S0_BY_M7
  `undef AXI_BV_S0_BY_M7
`endif 

`ifdef AXI_BV_S0_BY_M8
  `undef AXI_BV_S0_BY_M8
`endif 

`ifdef AXI_BV_S0_BY_M9
  `undef AXI_BV_S0_BY_M9
`endif 

`ifdef AXI_BV_S0_BY_M10
  `undef AXI_BV_S0_BY_M10
`endif 

`ifdef AXI_BV_S0_BY_M11
  `undef AXI_BV_S0_BY_M11
`endif 

`ifdef AXI_BV_S0_BY_M12
  `undef AXI_BV_S0_BY_M12
`endif 

`ifdef AXI_BV_S0_BY_M13
  `undef AXI_BV_S0_BY_M13
`endif 

`ifdef AXI_BV_S0_BY_M14
  `undef AXI_BV_S0_BY_M14
`endif 

`ifdef AXI_BV_S0_BY_M15
  `undef AXI_BV_S0_BY_M15
`endif 

`ifdef AXI_BV_S0_BY_M16
  `undef AXI_BV_S0_BY_M16
`endif 

`ifdef AXI_BV_S1_BY_M1
  `undef AXI_BV_S1_BY_M1
`endif 

`ifdef AXI_BV_S1_BY_M2
  `undef AXI_BV_S1_BY_M2
`endif 

`ifdef AXI_BV_S1_BY_M3
  `undef AXI_BV_S1_BY_M3
`endif 

`ifdef AXI_BV_S1_BY_M4
  `undef AXI_BV_S1_BY_M4
`endif 

`ifdef AXI_BV_S1_BY_M5
  `undef AXI_BV_S1_BY_M5
`endif 

`ifdef AXI_BV_S1_BY_M6
  `undef AXI_BV_S1_BY_M6
`endif 

`ifdef AXI_BV_S1_BY_M7
  `undef AXI_BV_S1_BY_M7
`endif 

`ifdef AXI_BV_S1_BY_M8
  `undef AXI_BV_S1_BY_M8
`endif 

`ifdef AXI_BV_S1_BY_M9
  `undef AXI_BV_S1_BY_M9
`endif 

`ifdef AXI_BV_S1_BY_M10
  `undef AXI_BV_S1_BY_M10
`endif 

`ifdef AXI_BV_S1_BY_M11
  `undef AXI_BV_S1_BY_M11
`endif 

`ifdef AXI_BV_S1_BY_M12
  `undef AXI_BV_S1_BY_M12
`endif 

`ifdef AXI_BV_S1_BY_M13
  `undef AXI_BV_S1_BY_M13
`endif 

`ifdef AXI_BV_S1_BY_M14
  `undef AXI_BV_S1_BY_M14
`endif 

`ifdef AXI_BV_S1_BY_M15
  `undef AXI_BV_S1_BY_M15
`endif 

`ifdef AXI_BV_S1_BY_M16
  `undef AXI_BV_S1_BY_M16
`endif 

`ifdef AXI_BV_S2_BY_M1
  `undef AXI_BV_S2_BY_M1
`endif 

`ifdef AXI_BV_S2_BY_M2
  `undef AXI_BV_S2_BY_M2
`endif 

`ifdef AXI_BV_S2_BY_M3
  `undef AXI_BV_S2_BY_M3
`endif 

`ifdef AXI_BV_S2_BY_M4
  `undef AXI_BV_S2_BY_M4
`endif 

`ifdef AXI_BV_S2_BY_M5
  `undef AXI_BV_S2_BY_M5
`endif 

`ifdef AXI_BV_S2_BY_M6
  `undef AXI_BV_S2_BY_M6
`endif 

`ifdef AXI_BV_S2_BY_M7
  `undef AXI_BV_S2_BY_M7
`endif 

`ifdef AXI_BV_S2_BY_M8
  `undef AXI_BV_S2_BY_M8
`endif 

`ifdef AXI_BV_S2_BY_M9
  `undef AXI_BV_S2_BY_M9
`endif 

`ifdef AXI_BV_S2_BY_M10
  `undef AXI_BV_S2_BY_M10
`endif 

`ifdef AXI_BV_S2_BY_M11
  `undef AXI_BV_S2_BY_M11
`endif 

`ifdef AXI_BV_S2_BY_M12
  `undef AXI_BV_S2_BY_M12
`endif 

`ifdef AXI_BV_S2_BY_M13
  `undef AXI_BV_S2_BY_M13
`endif 

`ifdef AXI_BV_S2_BY_M14
  `undef AXI_BV_S2_BY_M14
`endif 

`ifdef AXI_BV_S2_BY_M15
  `undef AXI_BV_S2_BY_M15
`endif 

`ifdef AXI_BV_S2_BY_M16
  `undef AXI_BV_S2_BY_M16
`endif 

`ifdef AXI_BV_S3_BY_M1
  `undef AXI_BV_S3_BY_M1
`endif 

`ifdef AXI_BV_S3_BY_M2
  `undef AXI_BV_S3_BY_M2
`endif 

`ifdef AXI_BV_S3_BY_M3
  `undef AXI_BV_S3_BY_M3
`endif 

`ifdef AXI_BV_S3_BY_M4
  `undef AXI_BV_S3_BY_M4
`endif 

`ifdef AXI_BV_S3_BY_M5
  `undef AXI_BV_S3_BY_M5
`endif 

`ifdef AXI_BV_S3_BY_M6
  `undef AXI_BV_S3_BY_M6
`endif 

`ifdef AXI_BV_S3_BY_M7
  `undef AXI_BV_S3_BY_M7
`endif 

`ifdef AXI_BV_S3_BY_M8
  `undef AXI_BV_S3_BY_M8
`endif 

`ifdef AXI_BV_S3_BY_M9
  `undef AXI_BV_S3_BY_M9
`endif 

`ifdef AXI_BV_S3_BY_M10
  `undef AXI_BV_S3_BY_M10
`endif 

`ifdef AXI_BV_S3_BY_M11
  `undef AXI_BV_S3_BY_M11
`endif 

`ifdef AXI_BV_S3_BY_M12
  `undef AXI_BV_S3_BY_M12
`endif 

`ifdef AXI_BV_S3_BY_M13
  `undef AXI_BV_S3_BY_M13
`endif 

`ifdef AXI_BV_S3_BY_M14
  `undef AXI_BV_S3_BY_M14
`endif 

`ifdef AXI_BV_S3_BY_M15
  `undef AXI_BV_S3_BY_M15
`endif 

`ifdef AXI_BV_S3_BY_M16
  `undef AXI_BV_S3_BY_M16
`endif 

`ifdef AXI_BV_S4_BY_M1
  `undef AXI_BV_S4_BY_M1
`endif 

`ifdef AXI_BV_S4_BY_M2
  `undef AXI_BV_S4_BY_M2
`endif 

`ifdef AXI_BV_S4_BY_M3
  `undef AXI_BV_S4_BY_M3
`endif 

`ifdef AXI_BV_S4_BY_M4
  `undef AXI_BV_S4_BY_M4
`endif 

`ifdef AXI_BV_S4_BY_M5
  `undef AXI_BV_S4_BY_M5
`endif 

`ifdef AXI_BV_S4_BY_M6
  `undef AXI_BV_S4_BY_M6
`endif 

`ifdef AXI_BV_S4_BY_M7
  `undef AXI_BV_S4_BY_M7
`endif 

`ifdef AXI_BV_S4_BY_M8
  `undef AXI_BV_S4_BY_M8
`endif 

`ifdef AXI_BV_S4_BY_M9
  `undef AXI_BV_S4_BY_M9
`endif 

`ifdef AXI_BV_S4_BY_M10
  `undef AXI_BV_S4_BY_M10
`endif 

`ifdef AXI_BV_S4_BY_M11
  `undef AXI_BV_S4_BY_M11
`endif 

`ifdef AXI_BV_S4_BY_M12
  `undef AXI_BV_S4_BY_M12
`endif 

`ifdef AXI_BV_S4_BY_M13
  `undef AXI_BV_S4_BY_M13
`endif 

`ifdef AXI_BV_S4_BY_M14
  `undef AXI_BV_S4_BY_M14
`endif 

`ifdef AXI_BV_S4_BY_M15
  `undef AXI_BV_S4_BY_M15
`endif 

`ifdef AXI_BV_S4_BY_M16
  `undef AXI_BV_S4_BY_M16
`endif 

`ifdef AXI_BV_S5_BY_M1
  `undef AXI_BV_S5_BY_M1
`endif 

`ifdef AXI_BV_S5_BY_M2
  `undef AXI_BV_S5_BY_M2
`endif 

`ifdef AXI_BV_S5_BY_M3
  `undef AXI_BV_S5_BY_M3
`endif 

`ifdef AXI_BV_S5_BY_M4
  `undef AXI_BV_S5_BY_M4
`endif 

`ifdef AXI_BV_S5_BY_M5
  `undef AXI_BV_S5_BY_M5
`endif 

`ifdef AXI_BV_S5_BY_M6
  `undef AXI_BV_S5_BY_M6
`endif 

`ifdef AXI_BV_S5_BY_M7
  `undef AXI_BV_S5_BY_M7
`endif 

`ifdef AXI_BV_S5_BY_M8
  `undef AXI_BV_S5_BY_M8
`endif 

`ifdef AXI_BV_S5_BY_M9
  `undef AXI_BV_S5_BY_M9
`endif 

`ifdef AXI_BV_S5_BY_M10
  `undef AXI_BV_S5_BY_M10
`endif 

`ifdef AXI_BV_S5_BY_M11
  `undef AXI_BV_S5_BY_M11
`endif 

`ifdef AXI_BV_S5_BY_M12
  `undef AXI_BV_S5_BY_M12
`endif 

`ifdef AXI_BV_S5_BY_M13
  `undef AXI_BV_S5_BY_M13
`endif 

`ifdef AXI_BV_S5_BY_M14
  `undef AXI_BV_S5_BY_M14
`endif 

`ifdef AXI_BV_S5_BY_M15
  `undef AXI_BV_S5_BY_M15
`endif 

`ifdef AXI_BV_S5_BY_M16
  `undef AXI_BV_S5_BY_M16
`endif 

`ifdef AXI_BV_S6_BY_M1
  `undef AXI_BV_S6_BY_M1
`endif 

`ifdef AXI_BV_S6_BY_M2
  `undef AXI_BV_S6_BY_M2
`endif 

`ifdef AXI_BV_S6_BY_M3
  `undef AXI_BV_S6_BY_M3
`endif 

`ifdef AXI_BV_S6_BY_M4
  `undef AXI_BV_S6_BY_M4
`endif 

`ifdef AXI_BV_S6_BY_M5
  `undef AXI_BV_S6_BY_M5
`endif 

`ifdef AXI_BV_S6_BY_M6
  `undef AXI_BV_S6_BY_M6
`endif 

`ifdef AXI_BV_S6_BY_M7
  `undef AXI_BV_S6_BY_M7
`endif 

`ifdef AXI_BV_S6_BY_M8
  `undef AXI_BV_S6_BY_M8
`endif 

`ifdef AXI_BV_S6_BY_M9
  `undef AXI_BV_S6_BY_M9
`endif 

`ifdef AXI_BV_S6_BY_M10
  `undef AXI_BV_S6_BY_M10
`endif 

`ifdef AXI_BV_S6_BY_M11
  `undef AXI_BV_S6_BY_M11
`endif 

`ifdef AXI_BV_S6_BY_M12
  `undef AXI_BV_S6_BY_M12
`endif 

`ifdef AXI_BV_S6_BY_M13
  `undef AXI_BV_S6_BY_M13
`endif 

`ifdef AXI_BV_S6_BY_M14
  `undef AXI_BV_S6_BY_M14
`endif 

`ifdef AXI_BV_S6_BY_M15
  `undef AXI_BV_S6_BY_M15
`endif 

`ifdef AXI_BV_S6_BY_M16
  `undef AXI_BV_S6_BY_M16
`endif 

`ifdef AXI_BV_S7_BY_M1
  `undef AXI_BV_S7_BY_M1
`endif 

`ifdef AXI_BV_S7_BY_M2
  `undef AXI_BV_S7_BY_M2
`endif 

`ifdef AXI_BV_S7_BY_M3
  `undef AXI_BV_S7_BY_M3
`endif 

`ifdef AXI_BV_S7_BY_M4
  `undef AXI_BV_S7_BY_M4
`endif 

`ifdef AXI_BV_S7_BY_M5
  `undef AXI_BV_S7_BY_M5
`endif 

`ifdef AXI_BV_S7_BY_M6
  `undef AXI_BV_S7_BY_M6
`endif 

`ifdef AXI_BV_S7_BY_M7
  `undef AXI_BV_S7_BY_M7
`endif 

`ifdef AXI_BV_S7_BY_M8
  `undef AXI_BV_S7_BY_M8
`endif 

`ifdef AXI_BV_S7_BY_M9
  `undef AXI_BV_S7_BY_M9
`endif 

`ifdef AXI_BV_S7_BY_M10
  `undef AXI_BV_S7_BY_M10
`endif 

`ifdef AXI_BV_S7_BY_M11
  `undef AXI_BV_S7_BY_M11
`endif 

`ifdef AXI_BV_S7_BY_M12
  `undef AXI_BV_S7_BY_M12
`endif 

`ifdef AXI_BV_S7_BY_M13
  `undef AXI_BV_S7_BY_M13
`endif 

`ifdef AXI_BV_S7_BY_M14
  `undef AXI_BV_S7_BY_M14
`endif 

`ifdef AXI_BV_S7_BY_M15
  `undef AXI_BV_S7_BY_M15
`endif 

`ifdef AXI_BV_S7_BY_M16
  `undef AXI_BV_S7_BY_M16
`endif 

`ifdef AXI_BV_S8_BY_M1
  `undef AXI_BV_S8_BY_M1
`endif 

`ifdef AXI_BV_S8_BY_M2
  `undef AXI_BV_S8_BY_M2
`endif 

`ifdef AXI_BV_S8_BY_M3
  `undef AXI_BV_S8_BY_M3
`endif 

`ifdef AXI_BV_S8_BY_M4
  `undef AXI_BV_S8_BY_M4
`endif 

`ifdef AXI_BV_S8_BY_M5
  `undef AXI_BV_S8_BY_M5
`endif 

`ifdef AXI_BV_S8_BY_M6
  `undef AXI_BV_S8_BY_M6
`endif 

`ifdef AXI_BV_S8_BY_M7
  `undef AXI_BV_S8_BY_M7
`endif 

`ifdef AXI_BV_S8_BY_M8
  `undef AXI_BV_S8_BY_M8
`endif 

`ifdef AXI_BV_S8_BY_M9
  `undef AXI_BV_S8_BY_M9
`endif 

`ifdef AXI_BV_S8_BY_M10
  `undef AXI_BV_S8_BY_M10
`endif 

`ifdef AXI_BV_S8_BY_M11
  `undef AXI_BV_S8_BY_M11
`endif 

`ifdef AXI_BV_S8_BY_M12
  `undef AXI_BV_S8_BY_M12
`endif 

`ifdef AXI_BV_S8_BY_M13
  `undef AXI_BV_S8_BY_M13
`endif 

`ifdef AXI_BV_S8_BY_M14
  `undef AXI_BV_S8_BY_M14
`endif 

`ifdef AXI_BV_S8_BY_M15
  `undef AXI_BV_S8_BY_M15
`endif 

`ifdef AXI_BV_S8_BY_M16
  `undef AXI_BV_S8_BY_M16
`endif 

`ifdef AXI_BV_S9_BY_M1
  `undef AXI_BV_S9_BY_M1
`endif 

`ifdef AXI_BV_S9_BY_M2
  `undef AXI_BV_S9_BY_M2
`endif 

`ifdef AXI_BV_S9_BY_M3
  `undef AXI_BV_S9_BY_M3
`endif 

`ifdef AXI_BV_S9_BY_M4
  `undef AXI_BV_S9_BY_M4
`endif 

`ifdef AXI_BV_S9_BY_M5
  `undef AXI_BV_S9_BY_M5
`endif 

`ifdef AXI_BV_S9_BY_M6
  `undef AXI_BV_S9_BY_M6
`endif 

`ifdef AXI_BV_S9_BY_M7
  `undef AXI_BV_S9_BY_M7
`endif 

`ifdef AXI_BV_S9_BY_M8
  `undef AXI_BV_S9_BY_M8
`endif 

`ifdef AXI_BV_S9_BY_M9
  `undef AXI_BV_S9_BY_M9
`endif 

`ifdef AXI_BV_S9_BY_M10
  `undef AXI_BV_S9_BY_M10
`endif 

`ifdef AXI_BV_S9_BY_M11
  `undef AXI_BV_S9_BY_M11
`endif 

`ifdef AXI_BV_S9_BY_M12
  `undef AXI_BV_S9_BY_M12
`endif 

`ifdef AXI_BV_S9_BY_M13
  `undef AXI_BV_S9_BY_M13
`endif 

`ifdef AXI_BV_S9_BY_M14
  `undef AXI_BV_S9_BY_M14
`endif 

`ifdef AXI_BV_S9_BY_M15
  `undef AXI_BV_S9_BY_M15
`endif 

`ifdef AXI_BV_S9_BY_M16
  `undef AXI_BV_S9_BY_M16
`endif 

`ifdef AXI_BV_S10_BY_M1
  `undef AXI_BV_S10_BY_M1
`endif 

`ifdef AXI_BV_S10_BY_M2
  `undef AXI_BV_S10_BY_M2
`endif 

`ifdef AXI_BV_S10_BY_M3
  `undef AXI_BV_S10_BY_M3
`endif 

`ifdef AXI_BV_S10_BY_M4
  `undef AXI_BV_S10_BY_M4
`endif 

`ifdef AXI_BV_S10_BY_M5
  `undef AXI_BV_S10_BY_M5
`endif 

`ifdef AXI_BV_S10_BY_M6
  `undef AXI_BV_S10_BY_M6
`endif 

`ifdef AXI_BV_S10_BY_M7
  `undef AXI_BV_S10_BY_M7
`endif 

`ifdef AXI_BV_S10_BY_M8
  `undef AXI_BV_S10_BY_M8
`endif 

`ifdef AXI_BV_S10_BY_M9
  `undef AXI_BV_S10_BY_M9
`endif 

`ifdef AXI_BV_S10_BY_M10
  `undef AXI_BV_S10_BY_M10
`endif 

`ifdef AXI_BV_S10_BY_M11
  `undef AXI_BV_S10_BY_M11
`endif 

`ifdef AXI_BV_S10_BY_M12
  `undef AXI_BV_S10_BY_M12
`endif 

`ifdef AXI_BV_S10_BY_M13
  `undef AXI_BV_S10_BY_M13
`endif 

`ifdef AXI_BV_S10_BY_M14
  `undef AXI_BV_S10_BY_M14
`endif 

`ifdef AXI_BV_S10_BY_M15
  `undef AXI_BV_S10_BY_M15
`endif 

`ifdef AXI_BV_S10_BY_M16
  `undef AXI_BV_S10_BY_M16
`endif 

`ifdef AXI_BV_S11_BY_M1
  `undef AXI_BV_S11_BY_M1
`endif 

`ifdef AXI_BV_S11_BY_M2
  `undef AXI_BV_S11_BY_M2
`endif 

`ifdef AXI_BV_S11_BY_M3
  `undef AXI_BV_S11_BY_M3
`endif 

`ifdef AXI_BV_S11_BY_M4
  `undef AXI_BV_S11_BY_M4
`endif 

`ifdef AXI_BV_S11_BY_M5
  `undef AXI_BV_S11_BY_M5
`endif 

`ifdef AXI_BV_S11_BY_M6
  `undef AXI_BV_S11_BY_M6
`endif 

`ifdef AXI_BV_S11_BY_M7
  `undef AXI_BV_S11_BY_M7
`endif 

`ifdef AXI_BV_S11_BY_M8
  `undef AXI_BV_S11_BY_M8
`endif 

`ifdef AXI_BV_S11_BY_M9
  `undef AXI_BV_S11_BY_M9
`endif 

`ifdef AXI_BV_S11_BY_M10
  `undef AXI_BV_S11_BY_M10
`endif 

`ifdef AXI_BV_S11_BY_M11
  `undef AXI_BV_S11_BY_M11
`endif 

`ifdef AXI_BV_S11_BY_M12
  `undef AXI_BV_S11_BY_M12
`endif 

`ifdef AXI_BV_S11_BY_M13
  `undef AXI_BV_S11_BY_M13
`endif 

`ifdef AXI_BV_S11_BY_M14
  `undef AXI_BV_S11_BY_M14
`endif 

`ifdef AXI_BV_S11_BY_M15
  `undef AXI_BV_S11_BY_M15
`endif 

`ifdef AXI_BV_S11_BY_M16
  `undef AXI_BV_S11_BY_M16
`endif 

`ifdef AXI_BV_S12_BY_M1
  `undef AXI_BV_S12_BY_M1
`endif 

`ifdef AXI_BV_S12_BY_M2
  `undef AXI_BV_S12_BY_M2
`endif 

`ifdef AXI_BV_S12_BY_M3
  `undef AXI_BV_S12_BY_M3
`endif 

`ifdef AXI_BV_S12_BY_M4
  `undef AXI_BV_S12_BY_M4
`endif 

`ifdef AXI_BV_S12_BY_M5
  `undef AXI_BV_S12_BY_M5
`endif 

`ifdef AXI_BV_S12_BY_M6
  `undef AXI_BV_S12_BY_M6
`endif 

`ifdef AXI_BV_S12_BY_M7
  `undef AXI_BV_S12_BY_M7
`endif 

`ifdef AXI_BV_S12_BY_M8
  `undef AXI_BV_S12_BY_M8
`endif 

`ifdef AXI_BV_S12_BY_M9
  `undef AXI_BV_S12_BY_M9
`endif 

`ifdef AXI_BV_S12_BY_M10
  `undef AXI_BV_S12_BY_M10
`endif 

`ifdef AXI_BV_S12_BY_M11
  `undef AXI_BV_S12_BY_M11
`endif 

`ifdef AXI_BV_S12_BY_M12
  `undef AXI_BV_S12_BY_M12
`endif 

`ifdef AXI_BV_S12_BY_M13
  `undef AXI_BV_S12_BY_M13
`endif 

`ifdef AXI_BV_S12_BY_M14
  `undef AXI_BV_S12_BY_M14
`endif 

`ifdef AXI_BV_S12_BY_M15
  `undef AXI_BV_S12_BY_M15
`endif 

`ifdef AXI_BV_S12_BY_M16
  `undef AXI_BV_S12_BY_M16
`endif 

`ifdef AXI_BV_S13_BY_M1
  `undef AXI_BV_S13_BY_M1
`endif 

`ifdef AXI_BV_S13_BY_M2
  `undef AXI_BV_S13_BY_M2
`endif 

`ifdef AXI_BV_S13_BY_M3
  `undef AXI_BV_S13_BY_M3
`endif 

`ifdef AXI_BV_S13_BY_M4
  `undef AXI_BV_S13_BY_M4
`endif 

`ifdef AXI_BV_S13_BY_M5
  `undef AXI_BV_S13_BY_M5
`endif 

`ifdef AXI_BV_S13_BY_M6
  `undef AXI_BV_S13_BY_M6
`endif 

`ifdef AXI_BV_S13_BY_M7
  `undef AXI_BV_S13_BY_M7
`endif 

`ifdef AXI_BV_S13_BY_M8
  `undef AXI_BV_S13_BY_M8
`endif 

`ifdef AXI_BV_S13_BY_M9
  `undef AXI_BV_S13_BY_M9
`endif 

`ifdef AXI_BV_S13_BY_M10
  `undef AXI_BV_S13_BY_M10
`endif 

`ifdef AXI_BV_S13_BY_M11
  `undef AXI_BV_S13_BY_M11
`endif 

`ifdef AXI_BV_S13_BY_M12
  `undef AXI_BV_S13_BY_M12
`endif 

`ifdef AXI_BV_S13_BY_M13
  `undef AXI_BV_S13_BY_M13
`endif 

`ifdef AXI_BV_S13_BY_M14
  `undef AXI_BV_S13_BY_M14
`endif 

`ifdef AXI_BV_S13_BY_M15
  `undef AXI_BV_S13_BY_M15
`endif 

`ifdef AXI_BV_S13_BY_M16
  `undef AXI_BV_S13_BY_M16
`endif 

`ifdef AXI_BV_S14_BY_M1
  `undef AXI_BV_S14_BY_M1
`endif 

`ifdef AXI_BV_S14_BY_M2
  `undef AXI_BV_S14_BY_M2
`endif 

`ifdef AXI_BV_S14_BY_M3
  `undef AXI_BV_S14_BY_M3
`endif 

`ifdef AXI_BV_S14_BY_M4
  `undef AXI_BV_S14_BY_M4
`endif 

`ifdef AXI_BV_S14_BY_M5
  `undef AXI_BV_S14_BY_M5
`endif 

`ifdef AXI_BV_S14_BY_M6
  `undef AXI_BV_S14_BY_M6
`endif 

`ifdef AXI_BV_S14_BY_M7
  `undef AXI_BV_S14_BY_M7
`endif 

`ifdef AXI_BV_S14_BY_M8
  `undef AXI_BV_S14_BY_M8
`endif 

`ifdef AXI_BV_S14_BY_M9
  `undef AXI_BV_S14_BY_M9
`endif 

`ifdef AXI_BV_S14_BY_M10
  `undef AXI_BV_S14_BY_M10
`endif 

`ifdef AXI_BV_S14_BY_M11
  `undef AXI_BV_S14_BY_M11
`endif 

`ifdef AXI_BV_S14_BY_M12
  `undef AXI_BV_S14_BY_M12
`endif 

`ifdef AXI_BV_S14_BY_M13
  `undef AXI_BV_S14_BY_M13
`endif 

`ifdef AXI_BV_S14_BY_M14
  `undef AXI_BV_S14_BY_M14
`endif 

`ifdef AXI_BV_S14_BY_M15
  `undef AXI_BV_S14_BY_M15
`endif 

`ifdef AXI_BV_S14_BY_M16
  `undef AXI_BV_S14_BY_M16
`endif 

`ifdef AXI_BV_S15_BY_M1
  `undef AXI_BV_S15_BY_M1
`endif 

`ifdef AXI_BV_S15_BY_M2
  `undef AXI_BV_S15_BY_M2
`endif 

`ifdef AXI_BV_S15_BY_M3
  `undef AXI_BV_S15_BY_M3
`endif 

`ifdef AXI_BV_S15_BY_M4
  `undef AXI_BV_S15_BY_M4
`endif 

`ifdef AXI_BV_S15_BY_M5
  `undef AXI_BV_S15_BY_M5
`endif 

`ifdef AXI_BV_S15_BY_M6
  `undef AXI_BV_S15_BY_M6
`endif 

`ifdef AXI_BV_S15_BY_M7
  `undef AXI_BV_S15_BY_M7
`endif 

`ifdef AXI_BV_S15_BY_M8
  `undef AXI_BV_S15_BY_M8
`endif 

`ifdef AXI_BV_S15_BY_M9
  `undef AXI_BV_S15_BY_M9
`endif 

`ifdef AXI_BV_S15_BY_M10
  `undef AXI_BV_S15_BY_M10
`endif 

`ifdef AXI_BV_S15_BY_M11
  `undef AXI_BV_S15_BY_M11
`endif 

`ifdef AXI_BV_S15_BY_M12
  `undef AXI_BV_S15_BY_M12
`endif 

`ifdef AXI_BV_S15_BY_M13
  `undef AXI_BV_S15_BY_M13
`endif 

`ifdef AXI_BV_S15_BY_M14
  `undef AXI_BV_S15_BY_M14
`endif 

`ifdef AXI_BV_S15_BY_M15
  `undef AXI_BV_S15_BY_M15
`endif 

`ifdef AXI_BV_S15_BY_M16
  `undef AXI_BV_S15_BY_M16
`endif 

`ifdef AXI_BV_S16_BY_M1
  `undef AXI_BV_S16_BY_M1
`endif 

`ifdef AXI_BV_S16_BY_M2
  `undef AXI_BV_S16_BY_M2
`endif 

`ifdef AXI_BV_S16_BY_M3
  `undef AXI_BV_S16_BY_M3
`endif 

`ifdef AXI_BV_S16_BY_M4
  `undef AXI_BV_S16_BY_M4
`endif 

`ifdef AXI_BV_S16_BY_M5
  `undef AXI_BV_S16_BY_M5
`endif 

`ifdef AXI_BV_S16_BY_M6
  `undef AXI_BV_S16_BY_M6
`endif 

`ifdef AXI_BV_S16_BY_M7
  `undef AXI_BV_S16_BY_M7
`endif 

`ifdef AXI_BV_S16_BY_M8
  `undef AXI_BV_S16_BY_M8
`endif 

`ifdef AXI_BV_S16_BY_M9
  `undef AXI_BV_S16_BY_M9
`endif 

`ifdef AXI_BV_S16_BY_M10
  `undef AXI_BV_S16_BY_M10
`endif 

`ifdef AXI_BV_S16_BY_M11
  `undef AXI_BV_S16_BY_M11
`endif 

`ifdef AXI_BV_S16_BY_M12
  `undef AXI_BV_S16_BY_M12
`endif 

`ifdef AXI_BV_S16_BY_M13
  `undef AXI_BV_S16_BY_M13
`endif 

`ifdef AXI_BV_S16_BY_M14
  `undef AXI_BV_S16_BY_M14
`endif 

`ifdef AXI_BV_S16_BY_M15
  `undef AXI_BV_S16_BY_M15
`endif 

`ifdef AXI_BV_S16_BY_M16
  `undef AXI_BV_S16_BY_M16
`endif 

`ifdef AXI_BV_S1_BY_ANY_M
  `undef AXI_BV_S1_BY_ANY_M
`endif 

`ifdef AXI_BV_S2_BY_ANY_M
  `undef AXI_BV_S2_BY_ANY_M
`endif 

`ifdef AXI_BV_S3_BY_ANY_M
  `undef AXI_BV_S3_BY_ANY_M
`endif 

`ifdef AXI_BV_S4_BY_ANY_M
  `undef AXI_BV_S4_BY_ANY_M
`endif 

`ifdef AXI_BV_S5_BY_ANY_M
  `undef AXI_BV_S5_BY_ANY_M
`endif 

`ifdef AXI_BV_S6_BY_ANY_M
  `undef AXI_BV_S6_BY_ANY_M
`endif 

`ifdef AXI_BV_S7_BY_ANY_M
  `undef AXI_BV_S7_BY_ANY_M
`endif 

`ifdef AXI_BV_S8_BY_ANY_M
  `undef AXI_BV_S8_BY_ANY_M
`endif 

`ifdef AXI_BV_S9_BY_ANY_M
  `undef AXI_BV_S9_BY_ANY_M
`endif 

`ifdef AXI_BV_S10_BY_ANY_M
  `undef AXI_BV_S10_BY_ANY_M
`endif 

`ifdef AXI_BV_S11_BY_ANY_M
  `undef AXI_BV_S11_BY_ANY_M
`endif 

`ifdef AXI_BV_S12_BY_ANY_M
  `undef AXI_BV_S12_BY_ANY_M
`endif 

`ifdef AXI_BV_S13_BY_ANY_M
  `undef AXI_BV_S13_BY_ANY_M
`endif 

`ifdef AXI_BV_S14_BY_ANY_M
  `undef AXI_BV_S14_BY_ANY_M
`endif 

`ifdef AXI_BV_S15_BY_ANY_M
  `undef AXI_BV_S15_BY_ANY_M
`endif 

`ifdef AXI_BV_S16_BY_ANY_M
  `undef AXI_BV_S16_BY_ANY_M
`endif 

`ifdef AXI_VV_S0_BY_M1
  `undef AXI_VV_S0_BY_M1
`endif 

`ifdef AXI_V_S0_BY_M1
  `undef AXI_V_S0_BY_M1
`endif 

`ifdef AXI_VV_S0_BY_M2
  `undef AXI_VV_S0_BY_M2
`endif 

`ifdef AXI_V_S0_BY_M2
  `undef AXI_V_S0_BY_M2
`endif 

`ifdef AXI_VV_S0_BY_M3
  `undef AXI_VV_S0_BY_M3
`endif 

`ifdef AXI_VV_S0_BY_M4
  `undef AXI_VV_S0_BY_M4
`endif 

`ifdef AXI_VV_S0_BY_M5
  `undef AXI_VV_S0_BY_M5
`endif 

`ifdef AXI_VV_S0_BY_M6
  `undef AXI_VV_S0_BY_M6
`endif 

`ifdef AXI_VV_S0_BY_M7
  `undef AXI_VV_S0_BY_M7
`endif 

`ifdef AXI_VV_S0_BY_M8
  `undef AXI_VV_S0_BY_M8
`endif 

`ifdef AXI_VV_S0_BY_M9
  `undef AXI_VV_S0_BY_M9
`endif 

`ifdef AXI_VV_S0_BY_M10
  `undef AXI_VV_S0_BY_M10
`endif 

`ifdef AXI_VV_S0_BY_M11
  `undef AXI_VV_S0_BY_M11
`endif 

`ifdef AXI_VV_S0_BY_M12
  `undef AXI_VV_S0_BY_M12
`endif 

`ifdef AXI_VV_S0_BY_M13
  `undef AXI_VV_S0_BY_M13
`endif 

`ifdef AXI_VV_S0_BY_M14
  `undef AXI_VV_S0_BY_M14
`endif 

`ifdef AXI_VV_S0_BY_M15
  `undef AXI_VV_S0_BY_M15
`endif 

`ifdef AXI_VV_S0_BY_M16
  `undef AXI_VV_S0_BY_M16
`endif 

`ifdef AXI_VV_S1_BY_M1
  `undef AXI_VV_S1_BY_M1
`endif 

`ifdef AXI_V_S1_BY_M1
  `undef AXI_V_S1_BY_M1
`endif 

`ifdef AXI_VV_S1_BY_M2
  `undef AXI_VV_S1_BY_M2
`endif 

`ifdef AXI_V_S1_BY_M2
  `undef AXI_V_S1_BY_M2
`endif 

`ifdef AXI_VV_S1_BY_M3
  `undef AXI_VV_S1_BY_M3
`endif 

`ifdef AXI_VV_S1_BY_M4
  `undef AXI_VV_S1_BY_M4
`endif 

`ifdef AXI_VV_S1_BY_M5
  `undef AXI_VV_S1_BY_M5
`endif 

`ifdef AXI_VV_S1_BY_M6
  `undef AXI_VV_S1_BY_M6
`endif 

`ifdef AXI_VV_S1_BY_M7
  `undef AXI_VV_S1_BY_M7
`endif 

`ifdef AXI_VV_S1_BY_M8
  `undef AXI_VV_S1_BY_M8
`endif 

`ifdef AXI_VV_S1_BY_M9
  `undef AXI_VV_S1_BY_M9
`endif 

`ifdef AXI_VV_S1_BY_M10
  `undef AXI_VV_S1_BY_M10
`endif 

`ifdef AXI_VV_S1_BY_M11
  `undef AXI_VV_S1_BY_M11
`endif 

`ifdef AXI_VV_S1_BY_M12
  `undef AXI_VV_S1_BY_M12
`endif 

`ifdef AXI_VV_S1_BY_M13
  `undef AXI_VV_S1_BY_M13
`endif 

`ifdef AXI_VV_S1_BY_M14
  `undef AXI_VV_S1_BY_M14
`endif 

`ifdef AXI_VV_S1_BY_M15
  `undef AXI_VV_S1_BY_M15
`endif 

`ifdef AXI_VV_S1_BY_M16
  `undef AXI_VV_S1_BY_M16
`endif 

`ifdef AXI_VV_S2_BY_M1
  `undef AXI_VV_S2_BY_M1
`endif 

`ifdef AXI_V_S2_BY_M1
  `undef AXI_V_S2_BY_M1
`endif 

`ifdef AXI_VV_S2_BY_M2
  `undef AXI_VV_S2_BY_M2
`endif 

`ifdef AXI_V_S2_BY_M2
  `undef AXI_V_S2_BY_M2
`endif 

`ifdef AXI_VV_S2_BY_M3
  `undef AXI_VV_S2_BY_M3
`endif 

`ifdef AXI_VV_S2_BY_M4
  `undef AXI_VV_S2_BY_M4
`endif 

`ifdef AXI_VV_S2_BY_M5
  `undef AXI_VV_S2_BY_M5
`endif 

`ifdef AXI_VV_S2_BY_M6
  `undef AXI_VV_S2_BY_M6
`endif 

`ifdef AXI_VV_S2_BY_M7
  `undef AXI_VV_S2_BY_M7
`endif 

`ifdef AXI_VV_S2_BY_M8
  `undef AXI_VV_S2_BY_M8
`endif 

`ifdef AXI_VV_S2_BY_M9
  `undef AXI_VV_S2_BY_M9
`endif 

`ifdef AXI_VV_S2_BY_M10
  `undef AXI_VV_S2_BY_M10
`endif 

`ifdef AXI_VV_S2_BY_M11
  `undef AXI_VV_S2_BY_M11
`endif 

`ifdef AXI_VV_S2_BY_M12
  `undef AXI_VV_S2_BY_M12
`endif 

`ifdef AXI_VV_S2_BY_M13
  `undef AXI_VV_S2_BY_M13
`endif 

`ifdef AXI_VV_S2_BY_M14
  `undef AXI_VV_S2_BY_M14
`endif 

`ifdef AXI_VV_S2_BY_M15
  `undef AXI_VV_S2_BY_M15
`endif 

`ifdef AXI_VV_S2_BY_M16
  `undef AXI_VV_S2_BY_M16
`endif 

`ifdef AXI_VV_S3_BY_M1
  `undef AXI_VV_S3_BY_M1
`endif 

`ifdef AXI_V_S3_BY_M1
  `undef AXI_V_S3_BY_M1
`endif 

`ifdef AXI_VV_S3_BY_M2
  `undef AXI_VV_S3_BY_M2
`endif 

`ifdef AXI_V_S3_BY_M2
  `undef AXI_V_S3_BY_M2
`endif 

`ifdef AXI_VV_S3_BY_M3
  `undef AXI_VV_S3_BY_M3
`endif 

`ifdef AXI_VV_S3_BY_M4
  `undef AXI_VV_S3_BY_M4
`endif 

`ifdef AXI_VV_S3_BY_M5
  `undef AXI_VV_S3_BY_M5
`endif 

`ifdef AXI_VV_S3_BY_M6
  `undef AXI_VV_S3_BY_M6
`endif 

`ifdef AXI_VV_S3_BY_M7
  `undef AXI_VV_S3_BY_M7
`endif 

`ifdef AXI_VV_S3_BY_M8
  `undef AXI_VV_S3_BY_M8
`endif 

`ifdef AXI_VV_S3_BY_M9
  `undef AXI_VV_S3_BY_M9
`endif 

`ifdef AXI_VV_S3_BY_M10
  `undef AXI_VV_S3_BY_M10
`endif 

`ifdef AXI_VV_S3_BY_M11
  `undef AXI_VV_S3_BY_M11
`endif 

`ifdef AXI_VV_S3_BY_M12
  `undef AXI_VV_S3_BY_M12
`endif 

`ifdef AXI_VV_S3_BY_M13
  `undef AXI_VV_S3_BY_M13
`endif 

`ifdef AXI_VV_S3_BY_M14
  `undef AXI_VV_S3_BY_M14
`endif 

`ifdef AXI_VV_S3_BY_M15
  `undef AXI_VV_S3_BY_M15
`endif 

`ifdef AXI_VV_S3_BY_M16
  `undef AXI_VV_S3_BY_M16
`endif 

`ifdef AXI_VV_S4_BY_M1
  `undef AXI_VV_S4_BY_M1
`endif 

`ifdef AXI_VV_S4_BY_M2
  `undef AXI_VV_S4_BY_M2
`endif 

`ifdef AXI_VV_S4_BY_M3
  `undef AXI_VV_S4_BY_M3
`endif 

`ifdef AXI_VV_S4_BY_M4
  `undef AXI_VV_S4_BY_M4
`endif 

`ifdef AXI_VV_S4_BY_M5
  `undef AXI_VV_S4_BY_M5
`endif 

`ifdef AXI_VV_S4_BY_M6
  `undef AXI_VV_S4_BY_M6
`endif 

`ifdef AXI_VV_S4_BY_M7
  `undef AXI_VV_S4_BY_M7
`endif 

`ifdef AXI_VV_S4_BY_M8
  `undef AXI_VV_S4_BY_M8
`endif 

`ifdef AXI_VV_S4_BY_M9
  `undef AXI_VV_S4_BY_M9
`endif 

`ifdef AXI_VV_S4_BY_M10
  `undef AXI_VV_S4_BY_M10
`endif 

`ifdef AXI_VV_S4_BY_M11
  `undef AXI_VV_S4_BY_M11
`endif 

`ifdef AXI_VV_S4_BY_M12
  `undef AXI_VV_S4_BY_M12
`endif 

`ifdef AXI_VV_S4_BY_M13
  `undef AXI_VV_S4_BY_M13
`endif 

`ifdef AXI_VV_S4_BY_M14
  `undef AXI_VV_S4_BY_M14
`endif 

`ifdef AXI_VV_S4_BY_M15
  `undef AXI_VV_S4_BY_M15
`endif 

`ifdef AXI_VV_S4_BY_M16
  `undef AXI_VV_S4_BY_M16
`endif 

`ifdef AXI_VV_S5_BY_M1
  `undef AXI_VV_S5_BY_M1
`endif 

`ifdef AXI_VV_S5_BY_M2
  `undef AXI_VV_S5_BY_M2
`endif 

`ifdef AXI_VV_S5_BY_M3
  `undef AXI_VV_S5_BY_M3
`endif 

`ifdef AXI_VV_S5_BY_M4
  `undef AXI_VV_S5_BY_M4
`endif 

`ifdef AXI_VV_S5_BY_M5
  `undef AXI_VV_S5_BY_M5
`endif 

`ifdef AXI_VV_S5_BY_M6
  `undef AXI_VV_S5_BY_M6
`endif 

`ifdef AXI_VV_S5_BY_M7
  `undef AXI_VV_S5_BY_M7
`endif 

`ifdef AXI_VV_S5_BY_M8
  `undef AXI_VV_S5_BY_M8
`endif 

`ifdef AXI_VV_S5_BY_M9
  `undef AXI_VV_S5_BY_M9
`endif 

`ifdef AXI_VV_S5_BY_M10
  `undef AXI_VV_S5_BY_M10
`endif 

`ifdef AXI_VV_S5_BY_M11
  `undef AXI_VV_S5_BY_M11
`endif 

`ifdef AXI_VV_S5_BY_M12
  `undef AXI_VV_S5_BY_M12
`endif 

`ifdef AXI_VV_S5_BY_M13
  `undef AXI_VV_S5_BY_M13
`endif 

`ifdef AXI_VV_S5_BY_M14
  `undef AXI_VV_S5_BY_M14
`endif 

`ifdef AXI_VV_S5_BY_M15
  `undef AXI_VV_S5_BY_M15
`endif 

`ifdef AXI_VV_S5_BY_M16
  `undef AXI_VV_S5_BY_M16
`endif 

`ifdef AXI_VV_S6_BY_M1
  `undef AXI_VV_S6_BY_M1
`endif 

`ifdef AXI_VV_S6_BY_M2
  `undef AXI_VV_S6_BY_M2
`endif 

`ifdef AXI_VV_S6_BY_M3
  `undef AXI_VV_S6_BY_M3
`endif 

`ifdef AXI_VV_S6_BY_M4
  `undef AXI_VV_S6_BY_M4
`endif 

`ifdef AXI_VV_S6_BY_M5
  `undef AXI_VV_S6_BY_M5
`endif 

`ifdef AXI_VV_S6_BY_M6
  `undef AXI_VV_S6_BY_M6
`endif 

`ifdef AXI_VV_S6_BY_M7
  `undef AXI_VV_S6_BY_M7
`endif 

`ifdef AXI_VV_S6_BY_M8
  `undef AXI_VV_S6_BY_M8
`endif 

`ifdef AXI_VV_S6_BY_M9
  `undef AXI_VV_S6_BY_M9
`endif 

`ifdef AXI_VV_S6_BY_M10
  `undef AXI_VV_S6_BY_M10
`endif 

`ifdef AXI_VV_S6_BY_M11
  `undef AXI_VV_S6_BY_M11
`endif 

`ifdef AXI_VV_S6_BY_M12
  `undef AXI_VV_S6_BY_M12
`endif 

`ifdef AXI_VV_S6_BY_M13
  `undef AXI_VV_S6_BY_M13
`endif 

`ifdef AXI_VV_S6_BY_M14
  `undef AXI_VV_S6_BY_M14
`endif 

`ifdef AXI_VV_S6_BY_M15
  `undef AXI_VV_S6_BY_M15
`endif 

`ifdef AXI_VV_S6_BY_M16
  `undef AXI_VV_S6_BY_M16
`endif 

`ifdef AXI_VV_S7_BY_M1
  `undef AXI_VV_S7_BY_M1
`endif 

`ifdef AXI_VV_S7_BY_M2
  `undef AXI_VV_S7_BY_M2
`endif 

`ifdef AXI_VV_S7_BY_M3
  `undef AXI_VV_S7_BY_M3
`endif 

`ifdef AXI_VV_S7_BY_M4
  `undef AXI_VV_S7_BY_M4
`endif 

`ifdef AXI_VV_S7_BY_M5
  `undef AXI_VV_S7_BY_M5
`endif 

`ifdef AXI_VV_S7_BY_M6
  `undef AXI_VV_S7_BY_M6
`endif 

`ifdef AXI_VV_S7_BY_M7
  `undef AXI_VV_S7_BY_M7
`endif 

`ifdef AXI_VV_S7_BY_M8
  `undef AXI_VV_S7_BY_M8
`endif 

`ifdef AXI_VV_S7_BY_M9
  `undef AXI_VV_S7_BY_M9
`endif 

`ifdef AXI_VV_S7_BY_M10
  `undef AXI_VV_S7_BY_M10
`endif 

`ifdef AXI_VV_S7_BY_M11
  `undef AXI_VV_S7_BY_M11
`endif 

`ifdef AXI_VV_S7_BY_M12
  `undef AXI_VV_S7_BY_M12
`endif 

`ifdef AXI_VV_S7_BY_M13
  `undef AXI_VV_S7_BY_M13
`endif 

`ifdef AXI_VV_S7_BY_M14
  `undef AXI_VV_S7_BY_M14
`endif 

`ifdef AXI_VV_S7_BY_M15
  `undef AXI_VV_S7_BY_M15
`endif 

`ifdef AXI_VV_S7_BY_M16
  `undef AXI_VV_S7_BY_M16
`endif 

`ifdef AXI_VV_S8_BY_M1
  `undef AXI_VV_S8_BY_M1
`endif 

`ifdef AXI_VV_S8_BY_M2
  `undef AXI_VV_S8_BY_M2
`endif 

`ifdef AXI_VV_S8_BY_M3
  `undef AXI_VV_S8_BY_M3
`endif 

`ifdef AXI_VV_S8_BY_M4
  `undef AXI_VV_S8_BY_M4
`endif 

`ifdef AXI_VV_S8_BY_M5
  `undef AXI_VV_S8_BY_M5
`endif 

`ifdef AXI_VV_S8_BY_M6
  `undef AXI_VV_S8_BY_M6
`endif 

`ifdef AXI_VV_S8_BY_M7
  `undef AXI_VV_S8_BY_M7
`endif 

`ifdef AXI_VV_S8_BY_M8
  `undef AXI_VV_S8_BY_M8
`endif 

`ifdef AXI_VV_S8_BY_M9
  `undef AXI_VV_S8_BY_M9
`endif 

`ifdef AXI_VV_S8_BY_M10
  `undef AXI_VV_S8_BY_M10
`endif 

`ifdef AXI_VV_S8_BY_M11
  `undef AXI_VV_S8_BY_M11
`endif 

`ifdef AXI_VV_S8_BY_M12
  `undef AXI_VV_S8_BY_M12
`endif 

`ifdef AXI_VV_S8_BY_M13
  `undef AXI_VV_S8_BY_M13
`endif 

`ifdef AXI_VV_S8_BY_M14
  `undef AXI_VV_S8_BY_M14
`endif 

`ifdef AXI_VV_S8_BY_M15
  `undef AXI_VV_S8_BY_M15
`endif 

`ifdef AXI_VV_S8_BY_M16
  `undef AXI_VV_S8_BY_M16
`endif 

`ifdef AXI_VV_S9_BY_M1
  `undef AXI_VV_S9_BY_M1
`endif 

`ifdef AXI_VV_S9_BY_M2
  `undef AXI_VV_S9_BY_M2
`endif 

`ifdef AXI_VV_S9_BY_M3
  `undef AXI_VV_S9_BY_M3
`endif 

`ifdef AXI_VV_S9_BY_M4
  `undef AXI_VV_S9_BY_M4
`endif 

`ifdef AXI_VV_S9_BY_M5
  `undef AXI_VV_S9_BY_M5
`endif 

`ifdef AXI_VV_S9_BY_M6
  `undef AXI_VV_S9_BY_M6
`endif 

`ifdef AXI_VV_S9_BY_M7
  `undef AXI_VV_S9_BY_M7
`endif 

`ifdef AXI_VV_S9_BY_M8
  `undef AXI_VV_S9_BY_M8
`endif 

`ifdef AXI_VV_S9_BY_M9
  `undef AXI_VV_S9_BY_M9
`endif 

`ifdef AXI_VV_S9_BY_M10
  `undef AXI_VV_S9_BY_M10
`endif 

`ifdef AXI_VV_S9_BY_M11
  `undef AXI_VV_S9_BY_M11
`endif 

`ifdef AXI_VV_S9_BY_M12
  `undef AXI_VV_S9_BY_M12
`endif 

`ifdef AXI_VV_S9_BY_M13
  `undef AXI_VV_S9_BY_M13
`endif 

`ifdef AXI_VV_S9_BY_M14
  `undef AXI_VV_S9_BY_M14
`endif 

`ifdef AXI_VV_S9_BY_M15
  `undef AXI_VV_S9_BY_M15
`endif 

`ifdef AXI_VV_S9_BY_M16
  `undef AXI_VV_S9_BY_M16
`endif 

`ifdef AXI_VV_S10_BY_M1
  `undef AXI_VV_S10_BY_M1
`endif 

`ifdef AXI_VV_S10_BY_M2
  `undef AXI_VV_S10_BY_M2
`endif 

`ifdef AXI_VV_S10_BY_M3
  `undef AXI_VV_S10_BY_M3
`endif 

`ifdef AXI_VV_S10_BY_M4
  `undef AXI_VV_S10_BY_M4
`endif 

`ifdef AXI_VV_S10_BY_M5
  `undef AXI_VV_S10_BY_M5
`endif 

`ifdef AXI_VV_S10_BY_M6
  `undef AXI_VV_S10_BY_M6
`endif 

`ifdef AXI_VV_S10_BY_M7
  `undef AXI_VV_S10_BY_M7
`endif 

`ifdef AXI_VV_S10_BY_M8
  `undef AXI_VV_S10_BY_M8
`endif 

`ifdef AXI_VV_S10_BY_M9
  `undef AXI_VV_S10_BY_M9
`endif 

`ifdef AXI_VV_S10_BY_M10
  `undef AXI_VV_S10_BY_M10
`endif 

`ifdef AXI_VV_S10_BY_M11
  `undef AXI_VV_S10_BY_M11
`endif 

`ifdef AXI_VV_S10_BY_M12
  `undef AXI_VV_S10_BY_M12
`endif 

`ifdef AXI_VV_S10_BY_M13
  `undef AXI_VV_S10_BY_M13
`endif 

`ifdef AXI_VV_S10_BY_M14
  `undef AXI_VV_S10_BY_M14
`endif 

`ifdef AXI_VV_S10_BY_M15
  `undef AXI_VV_S10_BY_M15
`endif 

`ifdef AXI_VV_S10_BY_M16
  `undef AXI_VV_S10_BY_M16
`endif 

`ifdef AXI_VV_S11_BY_M1
  `undef AXI_VV_S11_BY_M1
`endif 

`ifdef AXI_VV_S11_BY_M2
  `undef AXI_VV_S11_BY_M2
`endif 

`ifdef AXI_VV_S11_BY_M3
  `undef AXI_VV_S11_BY_M3
`endif 

`ifdef AXI_VV_S11_BY_M4
  `undef AXI_VV_S11_BY_M4
`endif 

`ifdef AXI_VV_S11_BY_M5
  `undef AXI_VV_S11_BY_M5
`endif 

`ifdef AXI_VV_S11_BY_M6
  `undef AXI_VV_S11_BY_M6
`endif 

`ifdef AXI_VV_S11_BY_M7
  `undef AXI_VV_S11_BY_M7
`endif 

`ifdef AXI_VV_S11_BY_M8
  `undef AXI_VV_S11_BY_M8
`endif 

`ifdef AXI_VV_S11_BY_M9
  `undef AXI_VV_S11_BY_M9
`endif 

`ifdef AXI_VV_S11_BY_M10
  `undef AXI_VV_S11_BY_M10
`endif 

`ifdef AXI_VV_S11_BY_M11
  `undef AXI_VV_S11_BY_M11
`endif 

`ifdef AXI_VV_S11_BY_M12
  `undef AXI_VV_S11_BY_M12
`endif 

`ifdef AXI_VV_S11_BY_M13
  `undef AXI_VV_S11_BY_M13
`endif 

`ifdef AXI_VV_S11_BY_M14
  `undef AXI_VV_S11_BY_M14
`endif 

`ifdef AXI_VV_S11_BY_M15
  `undef AXI_VV_S11_BY_M15
`endif 

`ifdef AXI_VV_S11_BY_M16
  `undef AXI_VV_S11_BY_M16
`endif 

`ifdef AXI_VV_S12_BY_M1
  `undef AXI_VV_S12_BY_M1
`endif 

`ifdef AXI_VV_S12_BY_M2
  `undef AXI_VV_S12_BY_M2
`endif 

`ifdef AXI_VV_S12_BY_M3
  `undef AXI_VV_S12_BY_M3
`endif 

`ifdef AXI_VV_S12_BY_M4
  `undef AXI_VV_S12_BY_M4
`endif 

`ifdef AXI_VV_S12_BY_M5
  `undef AXI_VV_S12_BY_M5
`endif 

`ifdef AXI_VV_S12_BY_M6
  `undef AXI_VV_S12_BY_M6
`endif 

`ifdef AXI_VV_S12_BY_M7
  `undef AXI_VV_S12_BY_M7
`endif 

`ifdef AXI_VV_S12_BY_M8
  `undef AXI_VV_S12_BY_M8
`endif 

`ifdef AXI_VV_S12_BY_M9
  `undef AXI_VV_S12_BY_M9
`endif 

`ifdef AXI_VV_S12_BY_M10
  `undef AXI_VV_S12_BY_M10
`endif 

`ifdef AXI_VV_S12_BY_M11
  `undef AXI_VV_S12_BY_M11
`endif 

`ifdef AXI_VV_S12_BY_M12
  `undef AXI_VV_S12_BY_M12
`endif 

`ifdef AXI_VV_S12_BY_M13
  `undef AXI_VV_S12_BY_M13
`endif 

`ifdef AXI_VV_S12_BY_M14
  `undef AXI_VV_S12_BY_M14
`endif 

`ifdef AXI_VV_S12_BY_M15
  `undef AXI_VV_S12_BY_M15
`endif 

`ifdef AXI_VV_S12_BY_M16
  `undef AXI_VV_S12_BY_M16
`endif 

`ifdef AXI_VV_S13_BY_M1
  `undef AXI_VV_S13_BY_M1
`endif 

`ifdef AXI_VV_S13_BY_M2
  `undef AXI_VV_S13_BY_M2
`endif 

`ifdef AXI_VV_S13_BY_M3
  `undef AXI_VV_S13_BY_M3
`endif 

`ifdef AXI_VV_S13_BY_M4
  `undef AXI_VV_S13_BY_M4
`endif 

`ifdef AXI_VV_S13_BY_M5
  `undef AXI_VV_S13_BY_M5
`endif 

`ifdef AXI_VV_S13_BY_M6
  `undef AXI_VV_S13_BY_M6
`endif 

`ifdef AXI_VV_S13_BY_M7
  `undef AXI_VV_S13_BY_M7
`endif 

`ifdef AXI_VV_S13_BY_M8
  `undef AXI_VV_S13_BY_M8
`endif 

`ifdef AXI_VV_S13_BY_M9
  `undef AXI_VV_S13_BY_M9
`endif 

`ifdef AXI_VV_S13_BY_M10
  `undef AXI_VV_S13_BY_M10
`endif 

`ifdef AXI_VV_S13_BY_M11
  `undef AXI_VV_S13_BY_M11
`endif 

`ifdef AXI_VV_S13_BY_M12
  `undef AXI_VV_S13_BY_M12
`endif 

`ifdef AXI_VV_S13_BY_M13
  `undef AXI_VV_S13_BY_M13
`endif 

`ifdef AXI_VV_S13_BY_M14
  `undef AXI_VV_S13_BY_M14
`endif 

`ifdef AXI_VV_S13_BY_M15
  `undef AXI_VV_S13_BY_M15
`endif 

`ifdef AXI_VV_S13_BY_M16
  `undef AXI_VV_S13_BY_M16
`endif 

`ifdef AXI_VV_S14_BY_M1
  `undef AXI_VV_S14_BY_M1
`endif 

`ifdef AXI_VV_S14_BY_M2
  `undef AXI_VV_S14_BY_M2
`endif 

`ifdef AXI_VV_S14_BY_M3
  `undef AXI_VV_S14_BY_M3
`endif 

`ifdef AXI_VV_S14_BY_M4
  `undef AXI_VV_S14_BY_M4
`endif 

`ifdef AXI_VV_S14_BY_M5
  `undef AXI_VV_S14_BY_M5
`endif 

`ifdef AXI_VV_S14_BY_M6
  `undef AXI_VV_S14_BY_M6
`endif 

`ifdef AXI_VV_S14_BY_M7
  `undef AXI_VV_S14_BY_M7
`endif 

`ifdef AXI_VV_S14_BY_M8
  `undef AXI_VV_S14_BY_M8
`endif 

`ifdef AXI_VV_S14_BY_M9
  `undef AXI_VV_S14_BY_M9
`endif 

`ifdef AXI_VV_S14_BY_M10
  `undef AXI_VV_S14_BY_M10
`endif 

`ifdef AXI_VV_S14_BY_M11
  `undef AXI_VV_S14_BY_M11
`endif 

`ifdef AXI_VV_S14_BY_M12
  `undef AXI_VV_S14_BY_M12
`endif 

`ifdef AXI_VV_S14_BY_M13
  `undef AXI_VV_S14_BY_M13
`endif 

`ifdef AXI_VV_S14_BY_M14
  `undef AXI_VV_S14_BY_M14
`endif 

`ifdef AXI_VV_S14_BY_M15
  `undef AXI_VV_S14_BY_M15
`endif 

`ifdef AXI_VV_S14_BY_M16
  `undef AXI_VV_S14_BY_M16
`endif 

`ifdef AXI_VV_S15_BY_M1
  `undef AXI_VV_S15_BY_M1
`endif 

`ifdef AXI_VV_S15_BY_M2
  `undef AXI_VV_S15_BY_M2
`endif 

`ifdef AXI_VV_S15_BY_M3
  `undef AXI_VV_S15_BY_M3
`endif 

`ifdef AXI_VV_S15_BY_M4
  `undef AXI_VV_S15_BY_M4
`endif 

`ifdef AXI_VV_S15_BY_M5
  `undef AXI_VV_S15_BY_M5
`endif 

`ifdef AXI_VV_S15_BY_M6
  `undef AXI_VV_S15_BY_M6
`endif 

`ifdef AXI_VV_S15_BY_M7
  `undef AXI_VV_S15_BY_M7
`endif 

`ifdef AXI_VV_S15_BY_M8
  `undef AXI_VV_S15_BY_M8
`endif 

`ifdef AXI_VV_S15_BY_M9
  `undef AXI_VV_S15_BY_M9
`endif 

`ifdef AXI_VV_S15_BY_M10
  `undef AXI_VV_S15_BY_M10
`endif 

`ifdef AXI_VV_S15_BY_M11
  `undef AXI_VV_S15_BY_M11
`endif 

`ifdef AXI_VV_S15_BY_M12
  `undef AXI_VV_S15_BY_M12
`endif 

`ifdef AXI_VV_S15_BY_M13
  `undef AXI_VV_S15_BY_M13
`endif 

`ifdef AXI_VV_S15_BY_M14
  `undef AXI_VV_S15_BY_M14
`endif 

`ifdef AXI_VV_S15_BY_M15
  `undef AXI_VV_S15_BY_M15
`endif 

`ifdef AXI_VV_S15_BY_M16
  `undef AXI_VV_S15_BY_M16
`endif 

`ifdef AXI_VV_S16_BY_M1
  `undef AXI_VV_S16_BY_M1
`endif 

`ifdef AXI_VV_S16_BY_M2
  `undef AXI_VV_S16_BY_M2
`endif 

`ifdef AXI_VV_S16_BY_M3
  `undef AXI_VV_S16_BY_M3
`endif 

`ifdef AXI_VV_S16_BY_M4
  `undef AXI_VV_S16_BY_M4
`endif 

`ifdef AXI_VV_S16_BY_M5
  `undef AXI_VV_S16_BY_M5
`endif 

`ifdef AXI_VV_S16_BY_M6
  `undef AXI_VV_S16_BY_M6
`endif 

`ifdef AXI_VV_S16_BY_M7
  `undef AXI_VV_S16_BY_M7
`endif 

`ifdef AXI_VV_S16_BY_M8
  `undef AXI_VV_S16_BY_M8
`endif 

`ifdef AXI_VV_S16_BY_M9
  `undef AXI_VV_S16_BY_M9
`endif 

`ifdef AXI_VV_S16_BY_M10
  `undef AXI_VV_S16_BY_M10
`endif 

`ifdef AXI_VV_S16_BY_M11
  `undef AXI_VV_S16_BY_M11
`endif 

`ifdef AXI_VV_S16_BY_M12
  `undef AXI_VV_S16_BY_M12
`endif 

`ifdef AXI_VV_S16_BY_M13
  `undef AXI_VV_S16_BY_M13
`endif 

`ifdef AXI_VV_S16_BY_M14
  `undef AXI_VV_S16_BY_M14
`endif 

`ifdef AXI_VV_S16_BY_M15
  `undef AXI_VV_S16_BY_M15
`endif 

`ifdef AXI_VV_S16_BY_M16
  `undef AXI_VV_S16_BY_M16
`endif 

`ifdef AXI_NMV_S1
  `undef AXI_NMV_S1
`endif 

`ifdef AXI_LOG2_NMV_S1
  `undef AXI_LOG2_NMV_S1
`endif 

`ifdef AXI_LOG2_NMP1V_S1
  `undef AXI_LOG2_NMP1V_S1
`endif 

`ifdef AXI_NMV_S2
  `undef AXI_NMV_S2
`endif 

`ifdef AXI_LOG2_NMV_S2
  `undef AXI_LOG2_NMV_S2
`endif 

`ifdef AXI_LOG2_NMP1V_S2
  `undef AXI_LOG2_NMP1V_S2
`endif 

`ifdef AXI_NMV_S3
  `undef AXI_NMV_S3
`endif 

`ifdef AXI_LOG2_NMV_S3
  `undef AXI_LOG2_NMV_S3
`endif 

`ifdef AXI_LOG2_NMP1V_S3
  `undef AXI_LOG2_NMP1V_S3
`endif 

`ifdef AXI_NMV_S4
  `undef AXI_NMV_S4
`endif 

`ifdef AXI_LOG2_NMV_S4
  `undef AXI_LOG2_NMV_S4
`endif 

`ifdef AXI_LOG2_NMP1V_S4
  `undef AXI_LOG2_NMP1V_S4
`endif 

`ifdef AXI_NMV_S5
  `undef AXI_NMV_S5
`endif 

`ifdef AXI_LOG2_NMV_S5
  `undef AXI_LOG2_NMV_S5
`endif 

`ifdef AXI_LOG2_NMP1V_S5
  `undef AXI_LOG2_NMP1V_S5
`endif 

`ifdef AXI_NMV_S6
  `undef AXI_NMV_S6
`endif 

`ifdef AXI_LOG2_NMV_S6
  `undef AXI_LOG2_NMV_S6
`endif 

`ifdef AXI_LOG2_NMP1V_S6
  `undef AXI_LOG2_NMP1V_S6
`endif 

`ifdef AXI_NMV_S7
  `undef AXI_NMV_S7
`endif 

`ifdef AXI_LOG2_NMV_S7
  `undef AXI_LOG2_NMV_S7
`endif 

`ifdef AXI_LOG2_NMP1V_S7
  `undef AXI_LOG2_NMP1V_S7
`endif 

`ifdef AXI_NMV_S8
  `undef AXI_NMV_S8
`endif 

`ifdef AXI_LOG2_NMV_S8
  `undef AXI_LOG2_NMV_S8
`endif 

`ifdef AXI_LOG2_NMP1V_S8
  `undef AXI_LOG2_NMP1V_S8
`endif 

`ifdef AXI_NMV_S9
  `undef AXI_NMV_S9
`endif 

`ifdef AXI_LOG2_NMV_S9
  `undef AXI_LOG2_NMV_S9
`endif 

`ifdef AXI_LOG2_NMP1V_S9
  `undef AXI_LOG2_NMP1V_S9
`endif 

`ifdef AXI_NMV_S10
  `undef AXI_NMV_S10
`endif 

`ifdef AXI_LOG2_NMV_S10
  `undef AXI_LOG2_NMV_S10
`endif 

`ifdef AXI_LOG2_NMP1V_S10
  `undef AXI_LOG2_NMP1V_S10
`endif 

`ifdef AXI_NMV_S11
  `undef AXI_NMV_S11
`endif 

`ifdef AXI_LOG2_NMV_S11
  `undef AXI_LOG2_NMV_S11
`endif 

`ifdef AXI_LOG2_NMP1V_S11
  `undef AXI_LOG2_NMP1V_S11
`endif 

`ifdef AXI_NMV_S12
  `undef AXI_NMV_S12
`endif 

`ifdef AXI_LOG2_NMV_S12
  `undef AXI_LOG2_NMV_S12
`endif 

`ifdef AXI_LOG2_NMP1V_S12
  `undef AXI_LOG2_NMP1V_S12
`endif 

`ifdef AXI_NMV_S13
  `undef AXI_NMV_S13
`endif 

`ifdef AXI_LOG2_NMV_S13
  `undef AXI_LOG2_NMV_S13
`endif 

`ifdef AXI_LOG2_NMP1V_S13
  `undef AXI_LOG2_NMP1V_S13
`endif 

`ifdef AXI_NMV_S14
  `undef AXI_NMV_S14
`endif 

`ifdef AXI_LOG2_NMV_S14
  `undef AXI_LOG2_NMV_S14
`endif 

`ifdef AXI_LOG2_NMP1V_S14
  `undef AXI_LOG2_NMP1V_S14
`endif 

`ifdef AXI_NMV_S15
  `undef AXI_NMV_S15
`endif 

`ifdef AXI_LOG2_NMV_S15
  `undef AXI_LOG2_NMV_S15
`endif 

`ifdef AXI_LOG2_NMP1V_S15
  `undef AXI_LOG2_NMP1V_S15
`endif 

`ifdef AXI_NMV_S16
  `undef AXI_NMV_S16
`endif 

`ifdef AXI_LOG2_NMV_S16
  `undef AXI_LOG2_NMV_S16
`endif 

`ifdef AXI_LOG2_NMP1V_S16
  `undef AXI_LOG2_NMP1V_S16
`endif 

`ifdef AXI_NSV_M1
  `undef AXI_NSV_M1
`endif 

`ifdef AXI_LOG2_NSV_M1
  `undef AXI_LOG2_NSV_M1
`endif 

`ifdef AXI_NSV_M2
  `undef AXI_NSV_M2
`endif 

`ifdef AXI_LOG2_NSV_M2
  `undef AXI_LOG2_NSV_M2
`endif 

`ifdef AXI_NSV_M3
  `undef AXI_NSV_M3
`endif 

`ifdef AXI_LOG2_NSV_M3
  `undef AXI_LOG2_NSV_M3
`endif 

`ifdef AXI_NSV_M4
  `undef AXI_NSV_M4
`endif 

`ifdef AXI_LOG2_NSV_M4
  `undef AXI_LOG2_NSV_M4
`endif 

`ifdef AXI_NSV_M5
  `undef AXI_NSV_M5
`endif 

`ifdef AXI_LOG2_NSV_M5
  `undef AXI_LOG2_NSV_M5
`endif 

`ifdef AXI_NSV_M6
  `undef AXI_NSV_M6
`endif 

`ifdef AXI_LOG2_NSV_M6
  `undef AXI_LOG2_NSV_M6
`endif 

`ifdef AXI_NSV_M7
  `undef AXI_NSV_M7
`endif 

`ifdef AXI_LOG2_NSV_M7
  `undef AXI_LOG2_NSV_M7
`endif 

`ifdef AXI_NSV_M8
  `undef AXI_NSV_M8
`endif 

`ifdef AXI_LOG2_NSV_M8
  `undef AXI_LOG2_NSV_M8
`endif 

`ifdef AXI_NSV_M9
  `undef AXI_NSV_M9
`endif 

`ifdef AXI_LOG2_NSV_M9
  `undef AXI_LOG2_NSV_M9
`endif 

`ifdef AXI_NSV_M10
  `undef AXI_NSV_M10
`endif 

`ifdef AXI_LOG2_NSV_M10
  `undef AXI_LOG2_NSV_M10
`endif 

`ifdef AXI_NSV_M11
  `undef AXI_NSV_M11
`endif 

`ifdef AXI_LOG2_NSV_M11
  `undef AXI_LOG2_NSV_M11
`endif 

`ifdef AXI_NSV_M12
  `undef AXI_NSV_M12
`endif 

`ifdef AXI_LOG2_NSV_M12
  `undef AXI_LOG2_NSV_M12
`endif 

`ifdef AXI_NSV_M13
  `undef AXI_NSV_M13
`endif 

`ifdef AXI_LOG2_NSV_M13
  `undef AXI_LOG2_NSV_M13
`endif 

`ifdef AXI_NSV_M14
  `undef AXI_NSV_M14
`endif 

`ifdef AXI_LOG2_NSV_M14
  `undef AXI_LOG2_NSV_M14
`endif 

`ifdef AXI_NSV_M15
  `undef AXI_NSV_M15
`endif 

`ifdef AXI_LOG2_NSV_M15
  `undef AXI_LOG2_NSV_M15
`endif 

`ifdef AXI_NSV_M16
  `undef AXI_NSV_M16
`endif 

`ifdef AXI_LOG2_NSV_M16
  `undef AXI_LOG2_NSV_M16
`endif 

`ifdef AXI_NNMV_S1
  `undef AXI_NNMV_S1
`endif 

`ifdef AXI_BNMV_S1
  `undef AXI_BNMV_S1
`endif 

`ifdef AXI_NNMV_S2
  `undef AXI_NNMV_S2
`endif 

`ifdef AXI_BNMV_S2
  `undef AXI_BNMV_S2
`endif 

`ifdef AXI_NNMV_S3
  `undef AXI_NNMV_S3
`endif 

`ifdef AXI_BNMV_S3
  `undef AXI_BNMV_S3
`endif 

`ifdef AXI_NNMV_S4
  `undef AXI_NNMV_S4
`endif 

`ifdef AXI_BNMV_S4
  `undef AXI_BNMV_S4
`endif 

`ifdef AXI_NNMV_S5
  `undef AXI_NNMV_S5
`endif 

`ifdef AXI_BNMV_S5
  `undef AXI_BNMV_S5
`endif 

`ifdef AXI_NNMV_S6
  `undef AXI_NNMV_S6
`endif 

`ifdef AXI_BNMV_S6
  `undef AXI_BNMV_S6
`endif 

`ifdef AXI_NNMV_S7
  `undef AXI_NNMV_S7
`endif 

`ifdef AXI_BNMV_S7
  `undef AXI_BNMV_S7
`endif 

`ifdef AXI_NNMV_S8
  `undef AXI_NNMV_S8
`endif 

`ifdef AXI_BNMV_S8
  `undef AXI_BNMV_S8
`endif 

`ifdef AXI_NNMV_S9
  `undef AXI_NNMV_S9
`endif 

`ifdef AXI_BNMV_S9
  `undef AXI_BNMV_S9
`endif 

`ifdef AXI_NNMV_S10
  `undef AXI_NNMV_S10
`endif 

`ifdef AXI_BNMV_S10
  `undef AXI_BNMV_S10
`endif 

`ifdef AXI_NNMV_S11
  `undef AXI_NNMV_S11
`endif 

`ifdef AXI_BNMV_S11
  `undef AXI_BNMV_S11
`endif 

`ifdef AXI_NNMV_S12
  `undef AXI_NNMV_S12
`endif 

`ifdef AXI_BNMV_S12
  `undef AXI_BNMV_S12
`endif 

`ifdef AXI_NNMV_S13
  `undef AXI_NNMV_S13
`endif 

`ifdef AXI_BNMV_S13
  `undef AXI_BNMV_S13
`endif 

`ifdef AXI_NNMV_S14
  `undef AXI_NNMV_S14
`endif 

`ifdef AXI_BNMV_S14
  `undef AXI_BNMV_S14
`endif 

`ifdef AXI_NNMV_S15
  `undef AXI_NNMV_S15
`endif 

`ifdef AXI_BNMV_S15
  `undef AXI_BNMV_S15
`endif 

`ifdef AXI_NNMV_S16
  `undef AXI_NNMV_S16
`endif 

`ifdef AXI_BNMV_S16
  `undef AXI_BNMV_S16
`endif 

`ifdef AXI_NSP1V_M1
  `undef AXI_NSP1V_M1
`endif 

`ifdef AXI_LOG2_NSP1V_M1
  `undef AXI_LOG2_NSP1V_M1
`endif 

`ifdef AXI_LOG2_NSP2V_M1
  `undef AXI_LOG2_NSP2V_M1
`endif 

`ifdef AXI_NSP1V_M2
  `undef AXI_NSP1V_M2
`endif 

`ifdef AXI_LOG2_NSP1V_M2
  `undef AXI_LOG2_NSP1V_M2
`endif 

`ifdef AXI_LOG2_NSP2V_M2
  `undef AXI_LOG2_NSP2V_M2
`endif 

`ifdef AXI_NSP1V_M3
  `undef AXI_NSP1V_M3
`endif 

`ifdef AXI_LOG2_NSP1V_M3
  `undef AXI_LOG2_NSP1V_M3
`endif 

`ifdef AXI_LOG2_NSP2V_M3
  `undef AXI_LOG2_NSP2V_M3
`endif 

`ifdef AXI_NSP1V_M4
  `undef AXI_NSP1V_M4
`endif 

`ifdef AXI_LOG2_NSP1V_M4
  `undef AXI_LOG2_NSP1V_M4
`endif 

`ifdef AXI_LOG2_NSP2V_M4
  `undef AXI_LOG2_NSP2V_M4
`endif 

`ifdef AXI_NSP1V_M5
  `undef AXI_NSP1V_M5
`endif 

`ifdef AXI_LOG2_NSP1V_M5
  `undef AXI_LOG2_NSP1V_M5
`endif 

`ifdef AXI_LOG2_NSP2V_M5
  `undef AXI_LOG2_NSP2V_M5
`endif 

`ifdef AXI_NSP1V_M6
  `undef AXI_NSP1V_M6
`endif 

`ifdef AXI_LOG2_NSP1V_M6
  `undef AXI_LOG2_NSP1V_M6
`endif 

`ifdef AXI_LOG2_NSP2V_M6
  `undef AXI_LOG2_NSP2V_M6
`endif 

`ifdef AXI_NSP1V_M7
  `undef AXI_NSP1V_M7
`endif 

`ifdef AXI_LOG2_NSP1V_M7
  `undef AXI_LOG2_NSP1V_M7
`endif 

`ifdef AXI_LOG2_NSP2V_M7
  `undef AXI_LOG2_NSP2V_M7
`endif 

`ifdef AXI_NSP1V_M8
  `undef AXI_NSP1V_M8
`endif 

`ifdef AXI_LOG2_NSP1V_M8
  `undef AXI_LOG2_NSP1V_M8
`endif 

`ifdef AXI_LOG2_NSP2V_M8
  `undef AXI_LOG2_NSP2V_M8
`endif 

`ifdef AXI_NSP1V_M9
  `undef AXI_NSP1V_M9
`endif 

`ifdef AXI_LOG2_NSP1V_M9
  `undef AXI_LOG2_NSP1V_M9
`endif 

`ifdef AXI_LOG2_NSP2V_M9
  `undef AXI_LOG2_NSP2V_M9
`endif 

`ifdef AXI_NSP1V_M10
  `undef AXI_NSP1V_M10
`endif 

`ifdef AXI_LOG2_NSP1V_M10
  `undef AXI_LOG2_NSP1V_M10
`endif 

`ifdef AXI_LOG2_NSP2V_M10
  `undef AXI_LOG2_NSP2V_M10
`endif 

`ifdef AXI_NSP1V_M11
  `undef AXI_NSP1V_M11
`endif 

`ifdef AXI_LOG2_NSP1V_M11
  `undef AXI_LOG2_NSP1V_M11
`endif 

`ifdef AXI_LOG2_NSP2V_M11
  `undef AXI_LOG2_NSP2V_M11
`endif 

`ifdef AXI_NSP1V_M12
  `undef AXI_NSP1V_M12
`endif 

`ifdef AXI_LOG2_NSP1V_M12
  `undef AXI_LOG2_NSP1V_M12
`endif 

`ifdef AXI_LOG2_NSP2V_M12
  `undef AXI_LOG2_NSP2V_M12
`endif 

`ifdef AXI_NSP1V_M13
  `undef AXI_NSP1V_M13
`endif 

`ifdef AXI_LOG2_NSP1V_M13
  `undef AXI_LOG2_NSP1V_M13
`endif 

`ifdef AXI_LOG2_NSP2V_M13
  `undef AXI_LOG2_NSP2V_M13
`endif 

`ifdef AXI_NSP1V_M14
  `undef AXI_NSP1V_M14
`endif 

`ifdef AXI_LOG2_NSP1V_M14
  `undef AXI_LOG2_NSP1V_M14
`endif 

`ifdef AXI_LOG2_NSP2V_M14
  `undef AXI_LOG2_NSP2V_M14
`endif 

`ifdef AXI_NSP1V_M15
  `undef AXI_NSP1V_M15
`endif 

`ifdef AXI_LOG2_NSP1V_M15
  `undef AXI_LOG2_NSP1V_M15
`endif 

`ifdef AXI_LOG2_NSP2V_M15
  `undef AXI_LOG2_NSP2V_M15
`endif 

`ifdef AXI_NSP1V_M16
  `undef AXI_NSP1V_M16
`endif 

`ifdef AXI_LOG2_NSP1V_M16
  `undef AXI_LOG2_NSP1V_M16
`endif 

`ifdef AXI_LOG2_NSP2V_M16
  `undef AXI_LOG2_NSP2V_M16
`endif 

`ifdef AXI_ALL_AR_LAYER_SHARED
  `undef AXI_ALL_AR_LAYER_SHARED
`endif 

`ifdef AXI_AR_LAYER_S0_M1
  `undef AXI_AR_LAYER_S0_M1
`endif 

`ifdef AXI_AR_LAYER_S0_M2
  `undef AXI_AR_LAYER_S0_M2
`endif 

`ifdef AXI_AR_LAYER_S0_M3
  `undef AXI_AR_LAYER_S0_M3
`endif 

`ifdef AXI_AR_LAYER_S0_M4
  `undef AXI_AR_LAYER_S0_M4
`endif 

`ifdef AXI_AR_LAYER_S0_M5
  `undef AXI_AR_LAYER_S0_M5
`endif 

`ifdef AXI_AR_LAYER_S0_M6
  `undef AXI_AR_LAYER_S0_M6
`endif 

`ifdef AXI_AR_LAYER_S0_M7
  `undef AXI_AR_LAYER_S0_M7
`endif 

`ifdef AXI_AR_LAYER_S0_M8
  `undef AXI_AR_LAYER_S0_M8
`endif 

`ifdef AXI_AR_LAYER_S0_M9
  `undef AXI_AR_LAYER_S0_M9
`endif 

`ifdef AXI_AR_LAYER_S0_M10
  `undef AXI_AR_LAYER_S0_M10
`endif 

`ifdef AXI_AR_LAYER_S0_M11
  `undef AXI_AR_LAYER_S0_M11
`endif 

`ifdef AXI_AR_LAYER_S0_M12
  `undef AXI_AR_LAYER_S0_M12
`endif 

`ifdef AXI_AR_LAYER_S0_M13
  `undef AXI_AR_LAYER_S0_M13
`endif 

`ifdef AXI_AR_LAYER_S0_M14
  `undef AXI_AR_LAYER_S0_M14
`endif 

`ifdef AXI_AR_LAYER_S0_M15
  `undef AXI_AR_LAYER_S0_M15
`endif 

`ifdef AXI_AR_LAYER_S0_M16
  `undef AXI_AR_LAYER_S0_M16
`endif 

`ifdef AXI_ALL_AW_LAYER_SHARED
  `undef AXI_ALL_AW_LAYER_SHARED
`endif 

`ifdef AXI_AW_LAYER_S0_M1
  `undef AXI_AW_LAYER_S0_M1
`endif 

`ifdef AXI_AW_LAYER_S0_M2
  `undef AXI_AW_LAYER_S0_M2
`endif 

`ifdef AXI_AW_LAYER_S0_M3
  `undef AXI_AW_LAYER_S0_M3
`endif 

`ifdef AXI_AW_LAYER_S0_M4
  `undef AXI_AW_LAYER_S0_M4
`endif 

`ifdef AXI_AW_LAYER_S0_M5
  `undef AXI_AW_LAYER_S0_M5
`endif 

`ifdef AXI_AW_LAYER_S0_M6
  `undef AXI_AW_LAYER_S0_M6
`endif 

`ifdef AXI_AW_LAYER_S0_M7
  `undef AXI_AW_LAYER_S0_M7
`endif 

`ifdef AXI_AW_LAYER_S0_M8
  `undef AXI_AW_LAYER_S0_M8
`endif 

`ifdef AXI_AW_LAYER_S0_M9
  `undef AXI_AW_LAYER_S0_M9
`endif 

`ifdef AXI_AW_LAYER_S0_M10
  `undef AXI_AW_LAYER_S0_M10
`endif 

`ifdef AXI_AW_LAYER_S0_M11
  `undef AXI_AW_LAYER_S0_M11
`endif 

`ifdef AXI_AW_LAYER_S0_M12
  `undef AXI_AW_LAYER_S0_M12
`endif 

`ifdef AXI_AW_LAYER_S0_M13
  `undef AXI_AW_LAYER_S0_M13
`endif 

`ifdef AXI_AW_LAYER_S0_M14
  `undef AXI_AW_LAYER_S0_M14
`endif 

`ifdef AXI_AW_LAYER_S0_M15
  `undef AXI_AW_LAYER_S0_M15
`endif 

`ifdef AXI_AW_LAYER_S0_M16
  `undef AXI_AW_LAYER_S0_M16
`endif 

`ifdef AXI_ALL_W_LAYER_SHARED
  `undef AXI_ALL_W_LAYER_SHARED
`endif 

`ifdef AXI_W_LAYER_S0_M1
  `undef AXI_W_LAYER_S0_M1
`endif 

`ifdef AXI_W_LAYER_S0_M2
  `undef AXI_W_LAYER_S0_M2
`endif 

`ifdef AXI_W_LAYER_S0_M3
  `undef AXI_W_LAYER_S0_M3
`endif 

`ifdef AXI_W_LAYER_S0_M4
  `undef AXI_W_LAYER_S0_M4
`endif 

`ifdef AXI_W_LAYER_S0_M5
  `undef AXI_W_LAYER_S0_M5
`endif 

`ifdef AXI_W_LAYER_S0_M6
  `undef AXI_W_LAYER_S0_M6
`endif 

`ifdef AXI_W_LAYER_S0_M7
  `undef AXI_W_LAYER_S0_M7
`endif 

`ifdef AXI_W_LAYER_S0_M8
  `undef AXI_W_LAYER_S0_M8
`endif 

`ifdef AXI_W_LAYER_S0_M9
  `undef AXI_W_LAYER_S0_M9
`endif 

`ifdef AXI_W_LAYER_S0_M10
  `undef AXI_W_LAYER_S0_M10
`endif 

`ifdef AXI_W_LAYER_S0_M11
  `undef AXI_W_LAYER_S0_M11
`endif 

`ifdef AXI_W_LAYER_S0_M12
  `undef AXI_W_LAYER_S0_M12
`endif 

`ifdef AXI_W_LAYER_S0_M13
  `undef AXI_W_LAYER_S0_M13
`endif 

`ifdef AXI_W_LAYER_S0_M14
  `undef AXI_W_LAYER_S0_M14
`endif 

`ifdef AXI_W_LAYER_S0_M15
  `undef AXI_W_LAYER_S0_M15
`endif 

`ifdef AXI_W_LAYER_S0_M16
  `undef AXI_W_LAYER_S0_M16
`endif 

`ifdef AXI_AR_LAYER_S1_M1
  `undef AXI_AR_LAYER_S1_M1
`endif 

`ifdef AXI_AR_LAYER_S1_M2
  `undef AXI_AR_LAYER_S1_M2
`endif 

`ifdef AXI_AR_LAYER_S1_M3
  `undef AXI_AR_LAYER_S1_M3
`endif 

`ifdef AXI_AR_LAYER_S1_M4
  `undef AXI_AR_LAYER_S1_M4
`endif 

`ifdef AXI_AR_LAYER_S1_M5
  `undef AXI_AR_LAYER_S1_M5
`endif 

`ifdef AXI_AR_LAYER_S1_M6
  `undef AXI_AR_LAYER_S1_M6
`endif 

`ifdef AXI_AR_LAYER_S1_M7
  `undef AXI_AR_LAYER_S1_M7
`endif 

`ifdef AXI_AR_LAYER_S1_M8
  `undef AXI_AR_LAYER_S1_M8
`endif 

`ifdef AXI_AR_LAYER_S1_M9
  `undef AXI_AR_LAYER_S1_M9
`endif 

`ifdef AXI_AR_LAYER_S1_M10
  `undef AXI_AR_LAYER_S1_M10
`endif 

`ifdef AXI_AR_LAYER_S1_M11
  `undef AXI_AR_LAYER_S1_M11
`endif 

`ifdef AXI_AR_LAYER_S1_M12
  `undef AXI_AR_LAYER_S1_M12
`endif 

`ifdef AXI_AR_LAYER_S1_M13
  `undef AXI_AR_LAYER_S1_M13
`endif 

`ifdef AXI_AR_LAYER_S1_M14
  `undef AXI_AR_LAYER_S1_M14
`endif 

`ifdef AXI_AR_LAYER_S1_M15
  `undef AXI_AR_LAYER_S1_M15
`endif 

`ifdef AXI_AR_LAYER_S1_M16
  `undef AXI_AR_LAYER_S1_M16
`endif 

`ifdef AXI_AW_LAYER_S1_M1
  `undef AXI_AW_LAYER_S1_M1
`endif 

`ifdef AXI_AW_LAYER_S1_M2
  `undef AXI_AW_LAYER_S1_M2
`endif 

`ifdef AXI_AW_LAYER_S1_M3
  `undef AXI_AW_LAYER_S1_M3
`endif 

`ifdef AXI_AW_LAYER_S1_M4
  `undef AXI_AW_LAYER_S1_M4
`endif 

`ifdef AXI_AW_LAYER_S1_M5
  `undef AXI_AW_LAYER_S1_M5
`endif 

`ifdef AXI_AW_LAYER_S1_M6
  `undef AXI_AW_LAYER_S1_M6
`endif 

`ifdef AXI_AW_LAYER_S1_M7
  `undef AXI_AW_LAYER_S1_M7
`endif 

`ifdef AXI_AW_LAYER_S1_M8
  `undef AXI_AW_LAYER_S1_M8
`endif 

`ifdef AXI_AW_LAYER_S1_M9
  `undef AXI_AW_LAYER_S1_M9
`endif 

`ifdef AXI_AW_LAYER_S1_M10
  `undef AXI_AW_LAYER_S1_M10
`endif 

`ifdef AXI_AW_LAYER_S1_M11
  `undef AXI_AW_LAYER_S1_M11
`endif 

`ifdef AXI_AW_LAYER_S1_M12
  `undef AXI_AW_LAYER_S1_M12
`endif 

`ifdef AXI_AW_LAYER_S1_M13
  `undef AXI_AW_LAYER_S1_M13
`endif 

`ifdef AXI_AW_LAYER_S1_M14
  `undef AXI_AW_LAYER_S1_M14
`endif 

`ifdef AXI_AW_LAYER_S1_M15
  `undef AXI_AW_LAYER_S1_M15
`endif 

`ifdef AXI_AW_LAYER_S1_M16
  `undef AXI_AW_LAYER_S1_M16
`endif 

`ifdef AXI_W_LAYER_S1_M1
  `undef AXI_W_LAYER_S1_M1
`endif 

`ifdef AXI_W_LAYER_S1_M2
  `undef AXI_W_LAYER_S1_M2
`endif 

`ifdef AXI_W_LAYER_S1_M3
  `undef AXI_W_LAYER_S1_M3
`endif 

`ifdef AXI_W_LAYER_S1_M4
  `undef AXI_W_LAYER_S1_M4
`endif 

`ifdef AXI_W_LAYER_S1_M5
  `undef AXI_W_LAYER_S1_M5
`endif 

`ifdef AXI_W_LAYER_S1_M6
  `undef AXI_W_LAYER_S1_M6
`endif 

`ifdef AXI_W_LAYER_S1_M7
  `undef AXI_W_LAYER_S1_M7
`endif 

`ifdef AXI_W_LAYER_S1_M8
  `undef AXI_W_LAYER_S1_M8
`endif 

`ifdef AXI_W_LAYER_S1_M9
  `undef AXI_W_LAYER_S1_M9
`endif 

`ifdef AXI_W_LAYER_S1_M10
  `undef AXI_W_LAYER_S1_M10
`endif 

`ifdef AXI_W_LAYER_S1_M11
  `undef AXI_W_LAYER_S1_M11
`endif 

`ifdef AXI_W_LAYER_S1_M12
  `undef AXI_W_LAYER_S1_M12
`endif 

`ifdef AXI_W_LAYER_S1_M13
  `undef AXI_W_LAYER_S1_M13
`endif 

`ifdef AXI_W_LAYER_S1_M14
  `undef AXI_W_LAYER_S1_M14
`endif 

`ifdef AXI_W_LAYER_S1_M15
  `undef AXI_W_LAYER_S1_M15
`endif 

`ifdef AXI_W_LAYER_S1_M16
  `undef AXI_W_LAYER_S1_M16
`endif 

`ifdef AXI_AR_LAYER_S2_M1
  `undef AXI_AR_LAYER_S2_M1
`endif 

`ifdef AXI_AR_LAYER_S2_M2
  `undef AXI_AR_LAYER_S2_M2
`endif 

`ifdef AXI_AR_LAYER_S2_M3
  `undef AXI_AR_LAYER_S2_M3
`endif 

`ifdef AXI_AR_LAYER_S2_M4
  `undef AXI_AR_LAYER_S2_M4
`endif 

`ifdef AXI_AR_LAYER_S2_M5
  `undef AXI_AR_LAYER_S2_M5
`endif 

`ifdef AXI_AR_LAYER_S2_M6
  `undef AXI_AR_LAYER_S2_M6
`endif 

`ifdef AXI_AR_LAYER_S2_M7
  `undef AXI_AR_LAYER_S2_M7
`endif 

`ifdef AXI_AR_LAYER_S2_M8
  `undef AXI_AR_LAYER_S2_M8
`endif 

`ifdef AXI_AR_LAYER_S2_M9
  `undef AXI_AR_LAYER_S2_M9
`endif 

`ifdef AXI_AR_LAYER_S2_M10
  `undef AXI_AR_LAYER_S2_M10
`endif 

`ifdef AXI_AR_LAYER_S2_M11
  `undef AXI_AR_LAYER_S2_M11
`endif 

`ifdef AXI_AR_LAYER_S2_M12
  `undef AXI_AR_LAYER_S2_M12
`endif 

`ifdef AXI_AR_LAYER_S2_M13
  `undef AXI_AR_LAYER_S2_M13
`endif 

`ifdef AXI_AR_LAYER_S2_M14
  `undef AXI_AR_LAYER_S2_M14
`endif 

`ifdef AXI_AR_LAYER_S2_M15
  `undef AXI_AR_LAYER_S2_M15
`endif 

`ifdef AXI_AR_LAYER_S2_M16
  `undef AXI_AR_LAYER_S2_M16
`endif 

`ifdef AXI_AW_LAYER_S2_M1
  `undef AXI_AW_LAYER_S2_M1
`endif 

`ifdef AXI_AW_LAYER_S2_M2
  `undef AXI_AW_LAYER_S2_M2
`endif 

`ifdef AXI_AW_LAYER_S2_M3
  `undef AXI_AW_LAYER_S2_M3
`endif 

`ifdef AXI_AW_LAYER_S2_M4
  `undef AXI_AW_LAYER_S2_M4
`endif 

`ifdef AXI_AW_LAYER_S2_M5
  `undef AXI_AW_LAYER_S2_M5
`endif 

`ifdef AXI_AW_LAYER_S2_M6
  `undef AXI_AW_LAYER_S2_M6
`endif 

`ifdef AXI_AW_LAYER_S2_M7
  `undef AXI_AW_LAYER_S2_M7
`endif 

`ifdef AXI_AW_LAYER_S2_M8
  `undef AXI_AW_LAYER_S2_M8
`endif 

`ifdef AXI_AW_LAYER_S2_M9
  `undef AXI_AW_LAYER_S2_M9
`endif 

`ifdef AXI_AW_LAYER_S2_M10
  `undef AXI_AW_LAYER_S2_M10
`endif 

`ifdef AXI_AW_LAYER_S2_M11
  `undef AXI_AW_LAYER_S2_M11
`endif 

`ifdef AXI_AW_LAYER_S2_M12
  `undef AXI_AW_LAYER_S2_M12
`endif 

`ifdef AXI_AW_LAYER_S2_M13
  `undef AXI_AW_LAYER_S2_M13
`endif 

`ifdef AXI_AW_LAYER_S2_M14
  `undef AXI_AW_LAYER_S2_M14
`endif 

`ifdef AXI_AW_LAYER_S2_M15
  `undef AXI_AW_LAYER_S2_M15
`endif 

`ifdef AXI_AW_LAYER_S2_M16
  `undef AXI_AW_LAYER_S2_M16
`endif 

`ifdef AXI_W_LAYER_S2_M1
  `undef AXI_W_LAYER_S2_M1
`endif 

`ifdef AXI_W_LAYER_S2_M2
  `undef AXI_W_LAYER_S2_M2
`endif 

`ifdef AXI_W_LAYER_S2_M3
  `undef AXI_W_LAYER_S2_M3
`endif 

`ifdef AXI_W_LAYER_S2_M4
  `undef AXI_W_LAYER_S2_M4
`endif 

`ifdef AXI_W_LAYER_S2_M5
  `undef AXI_W_LAYER_S2_M5
`endif 

`ifdef AXI_W_LAYER_S2_M6
  `undef AXI_W_LAYER_S2_M6
`endif 

`ifdef AXI_W_LAYER_S2_M7
  `undef AXI_W_LAYER_S2_M7
`endif 

`ifdef AXI_W_LAYER_S2_M8
  `undef AXI_W_LAYER_S2_M8
`endif 

`ifdef AXI_W_LAYER_S2_M9
  `undef AXI_W_LAYER_S2_M9
`endif 

`ifdef AXI_W_LAYER_S2_M10
  `undef AXI_W_LAYER_S2_M10
`endif 

`ifdef AXI_W_LAYER_S2_M11
  `undef AXI_W_LAYER_S2_M11
`endif 

`ifdef AXI_W_LAYER_S2_M12
  `undef AXI_W_LAYER_S2_M12
`endif 

`ifdef AXI_W_LAYER_S2_M13
  `undef AXI_W_LAYER_S2_M13
`endif 

`ifdef AXI_W_LAYER_S2_M14
  `undef AXI_W_LAYER_S2_M14
`endif 

`ifdef AXI_W_LAYER_S2_M15
  `undef AXI_W_LAYER_S2_M15
`endif 

`ifdef AXI_W_LAYER_S2_M16
  `undef AXI_W_LAYER_S2_M16
`endif 

`ifdef AXI_AR_LAYER_S3_M1
  `undef AXI_AR_LAYER_S3_M1
`endif 

`ifdef AXI_AR_LAYER_S3_M2
  `undef AXI_AR_LAYER_S3_M2
`endif 

`ifdef AXI_AR_LAYER_S3_M3
  `undef AXI_AR_LAYER_S3_M3
`endif 

`ifdef AXI_AR_LAYER_S3_M4
  `undef AXI_AR_LAYER_S3_M4
`endif 

`ifdef AXI_AR_LAYER_S3_M5
  `undef AXI_AR_LAYER_S3_M5
`endif 

`ifdef AXI_AR_LAYER_S3_M6
  `undef AXI_AR_LAYER_S3_M6
`endif 

`ifdef AXI_AR_LAYER_S3_M7
  `undef AXI_AR_LAYER_S3_M7
`endif 

`ifdef AXI_AR_LAYER_S3_M8
  `undef AXI_AR_LAYER_S3_M8
`endif 

`ifdef AXI_AR_LAYER_S3_M9
  `undef AXI_AR_LAYER_S3_M9
`endif 

`ifdef AXI_AR_LAYER_S3_M10
  `undef AXI_AR_LAYER_S3_M10
`endif 

`ifdef AXI_AR_LAYER_S3_M11
  `undef AXI_AR_LAYER_S3_M11
`endif 

`ifdef AXI_AR_LAYER_S3_M12
  `undef AXI_AR_LAYER_S3_M12
`endif 

`ifdef AXI_AR_LAYER_S3_M13
  `undef AXI_AR_LAYER_S3_M13
`endif 

`ifdef AXI_AR_LAYER_S3_M14
  `undef AXI_AR_LAYER_S3_M14
`endif 

`ifdef AXI_AR_LAYER_S3_M15
  `undef AXI_AR_LAYER_S3_M15
`endif 

`ifdef AXI_AR_LAYER_S3_M16
  `undef AXI_AR_LAYER_S3_M16
`endif 

`ifdef AXI_AW_LAYER_S3_M1
  `undef AXI_AW_LAYER_S3_M1
`endif 

`ifdef AXI_AW_LAYER_S3_M2
  `undef AXI_AW_LAYER_S3_M2
`endif 

`ifdef AXI_AW_LAYER_S3_M3
  `undef AXI_AW_LAYER_S3_M3
`endif 

`ifdef AXI_AW_LAYER_S3_M4
  `undef AXI_AW_LAYER_S3_M4
`endif 

`ifdef AXI_AW_LAYER_S3_M5
  `undef AXI_AW_LAYER_S3_M5
`endif 

`ifdef AXI_AW_LAYER_S3_M6
  `undef AXI_AW_LAYER_S3_M6
`endif 

`ifdef AXI_AW_LAYER_S3_M7
  `undef AXI_AW_LAYER_S3_M7
`endif 

`ifdef AXI_AW_LAYER_S3_M8
  `undef AXI_AW_LAYER_S3_M8
`endif 

`ifdef AXI_AW_LAYER_S3_M9
  `undef AXI_AW_LAYER_S3_M9
`endif 

`ifdef AXI_AW_LAYER_S3_M10
  `undef AXI_AW_LAYER_S3_M10
`endif 

`ifdef AXI_AW_LAYER_S3_M11
  `undef AXI_AW_LAYER_S3_M11
`endif 

`ifdef AXI_AW_LAYER_S3_M12
  `undef AXI_AW_LAYER_S3_M12
`endif 

`ifdef AXI_AW_LAYER_S3_M13
  `undef AXI_AW_LAYER_S3_M13
`endif 

`ifdef AXI_AW_LAYER_S3_M14
  `undef AXI_AW_LAYER_S3_M14
`endif 

`ifdef AXI_AW_LAYER_S3_M15
  `undef AXI_AW_LAYER_S3_M15
`endif 

`ifdef AXI_AW_LAYER_S3_M16
  `undef AXI_AW_LAYER_S3_M16
`endif 

`ifdef AXI_W_LAYER_S3_M1
  `undef AXI_W_LAYER_S3_M1
`endif 

`ifdef AXI_W_LAYER_S3_M2
  `undef AXI_W_LAYER_S3_M2
`endif 

`ifdef AXI_W_LAYER_S3_M3
  `undef AXI_W_LAYER_S3_M3
`endif 

`ifdef AXI_W_LAYER_S3_M4
  `undef AXI_W_LAYER_S3_M4
`endif 

`ifdef AXI_W_LAYER_S3_M5
  `undef AXI_W_LAYER_S3_M5
`endif 

`ifdef AXI_W_LAYER_S3_M6
  `undef AXI_W_LAYER_S3_M6
`endif 

`ifdef AXI_W_LAYER_S3_M7
  `undef AXI_W_LAYER_S3_M7
`endif 

`ifdef AXI_W_LAYER_S3_M8
  `undef AXI_W_LAYER_S3_M8
`endif 

`ifdef AXI_W_LAYER_S3_M9
  `undef AXI_W_LAYER_S3_M9
`endif 

`ifdef AXI_W_LAYER_S3_M10
  `undef AXI_W_LAYER_S3_M10
`endif 

`ifdef AXI_W_LAYER_S3_M11
  `undef AXI_W_LAYER_S3_M11
`endif 

`ifdef AXI_W_LAYER_S3_M12
  `undef AXI_W_LAYER_S3_M12
`endif 

`ifdef AXI_W_LAYER_S3_M13
  `undef AXI_W_LAYER_S3_M13
`endif 

`ifdef AXI_W_LAYER_S3_M14
  `undef AXI_W_LAYER_S3_M14
`endif 

`ifdef AXI_W_LAYER_S3_M15
  `undef AXI_W_LAYER_S3_M15
`endif 

`ifdef AXI_W_LAYER_S3_M16
  `undef AXI_W_LAYER_S3_M16
`endif 

`ifdef AXI_AR_LAYER_S4_M1
  `undef AXI_AR_LAYER_S4_M1
`endif 

`ifdef AXI_AR_LAYER_S4_M2
  `undef AXI_AR_LAYER_S4_M2
`endif 

`ifdef AXI_AR_LAYER_S4_M3
  `undef AXI_AR_LAYER_S4_M3
`endif 

`ifdef AXI_AR_LAYER_S4_M4
  `undef AXI_AR_LAYER_S4_M4
`endif 

`ifdef AXI_AR_LAYER_S4_M5
  `undef AXI_AR_LAYER_S4_M5
`endif 

`ifdef AXI_AR_LAYER_S4_M6
  `undef AXI_AR_LAYER_S4_M6
`endif 

`ifdef AXI_AR_LAYER_S4_M7
  `undef AXI_AR_LAYER_S4_M7
`endif 

`ifdef AXI_AR_LAYER_S4_M8
  `undef AXI_AR_LAYER_S4_M8
`endif 

`ifdef AXI_AR_LAYER_S4_M9
  `undef AXI_AR_LAYER_S4_M9
`endif 

`ifdef AXI_AR_LAYER_S4_M10
  `undef AXI_AR_LAYER_S4_M10
`endif 

`ifdef AXI_AR_LAYER_S4_M11
  `undef AXI_AR_LAYER_S4_M11
`endif 

`ifdef AXI_AR_LAYER_S4_M12
  `undef AXI_AR_LAYER_S4_M12
`endif 

`ifdef AXI_AR_LAYER_S4_M13
  `undef AXI_AR_LAYER_S4_M13
`endif 

`ifdef AXI_AR_LAYER_S4_M14
  `undef AXI_AR_LAYER_S4_M14
`endif 

`ifdef AXI_AR_LAYER_S4_M15
  `undef AXI_AR_LAYER_S4_M15
`endif 

`ifdef AXI_AR_LAYER_S4_M16
  `undef AXI_AR_LAYER_S4_M16
`endif 

`ifdef AXI_AW_LAYER_S4_M1
  `undef AXI_AW_LAYER_S4_M1
`endif 

`ifdef AXI_AW_LAYER_S4_M2
  `undef AXI_AW_LAYER_S4_M2
`endif 

`ifdef AXI_AW_LAYER_S4_M3
  `undef AXI_AW_LAYER_S4_M3
`endif 

`ifdef AXI_AW_LAYER_S4_M4
  `undef AXI_AW_LAYER_S4_M4
`endif 

`ifdef AXI_AW_LAYER_S4_M5
  `undef AXI_AW_LAYER_S4_M5
`endif 

`ifdef AXI_AW_LAYER_S4_M6
  `undef AXI_AW_LAYER_S4_M6
`endif 

`ifdef AXI_AW_LAYER_S4_M7
  `undef AXI_AW_LAYER_S4_M7
`endif 

`ifdef AXI_AW_LAYER_S4_M8
  `undef AXI_AW_LAYER_S4_M8
`endif 

`ifdef AXI_AW_LAYER_S4_M9
  `undef AXI_AW_LAYER_S4_M9
`endif 

`ifdef AXI_AW_LAYER_S4_M10
  `undef AXI_AW_LAYER_S4_M10
`endif 

`ifdef AXI_AW_LAYER_S4_M11
  `undef AXI_AW_LAYER_S4_M11
`endif 

`ifdef AXI_AW_LAYER_S4_M12
  `undef AXI_AW_LAYER_S4_M12
`endif 

`ifdef AXI_AW_LAYER_S4_M13
  `undef AXI_AW_LAYER_S4_M13
`endif 

`ifdef AXI_AW_LAYER_S4_M14
  `undef AXI_AW_LAYER_S4_M14
`endif 

`ifdef AXI_AW_LAYER_S4_M15
  `undef AXI_AW_LAYER_S4_M15
`endif 

`ifdef AXI_AW_LAYER_S4_M16
  `undef AXI_AW_LAYER_S4_M16
`endif 

`ifdef AXI_W_LAYER_S4_M1
  `undef AXI_W_LAYER_S4_M1
`endif 

`ifdef AXI_W_LAYER_S4_M2
  `undef AXI_W_LAYER_S4_M2
`endif 

`ifdef AXI_W_LAYER_S4_M3
  `undef AXI_W_LAYER_S4_M3
`endif 

`ifdef AXI_W_LAYER_S4_M4
  `undef AXI_W_LAYER_S4_M4
`endif 

`ifdef AXI_W_LAYER_S4_M5
  `undef AXI_W_LAYER_S4_M5
`endif 

`ifdef AXI_W_LAYER_S4_M6
  `undef AXI_W_LAYER_S4_M6
`endif 

`ifdef AXI_W_LAYER_S4_M7
  `undef AXI_W_LAYER_S4_M7
`endif 

`ifdef AXI_W_LAYER_S4_M8
  `undef AXI_W_LAYER_S4_M8
`endif 

`ifdef AXI_W_LAYER_S4_M9
  `undef AXI_W_LAYER_S4_M9
`endif 

`ifdef AXI_W_LAYER_S4_M10
  `undef AXI_W_LAYER_S4_M10
`endif 

`ifdef AXI_W_LAYER_S4_M11
  `undef AXI_W_LAYER_S4_M11
`endif 

`ifdef AXI_W_LAYER_S4_M12
  `undef AXI_W_LAYER_S4_M12
`endif 

`ifdef AXI_W_LAYER_S4_M13
  `undef AXI_W_LAYER_S4_M13
`endif 

`ifdef AXI_W_LAYER_S4_M14
  `undef AXI_W_LAYER_S4_M14
`endif 

`ifdef AXI_W_LAYER_S4_M15
  `undef AXI_W_LAYER_S4_M15
`endif 

`ifdef AXI_W_LAYER_S4_M16
  `undef AXI_W_LAYER_S4_M16
`endif 

`ifdef AXI_AR_LAYER_S5_M1
  `undef AXI_AR_LAYER_S5_M1
`endif 

`ifdef AXI_AR_LAYER_S5_M2
  `undef AXI_AR_LAYER_S5_M2
`endif 

`ifdef AXI_AR_LAYER_S5_M3
  `undef AXI_AR_LAYER_S5_M3
`endif 

`ifdef AXI_AR_LAYER_S5_M4
  `undef AXI_AR_LAYER_S5_M4
`endif 

`ifdef AXI_AR_LAYER_S5_M5
  `undef AXI_AR_LAYER_S5_M5
`endif 

`ifdef AXI_AR_LAYER_S5_M6
  `undef AXI_AR_LAYER_S5_M6
`endif 

`ifdef AXI_AR_LAYER_S5_M7
  `undef AXI_AR_LAYER_S5_M7
`endif 

`ifdef AXI_AR_LAYER_S5_M8
  `undef AXI_AR_LAYER_S5_M8
`endif 

`ifdef AXI_AR_LAYER_S5_M9
  `undef AXI_AR_LAYER_S5_M9
`endif 

`ifdef AXI_AR_LAYER_S5_M10
  `undef AXI_AR_LAYER_S5_M10
`endif 

`ifdef AXI_AR_LAYER_S5_M11
  `undef AXI_AR_LAYER_S5_M11
`endif 

`ifdef AXI_AR_LAYER_S5_M12
  `undef AXI_AR_LAYER_S5_M12
`endif 

`ifdef AXI_AR_LAYER_S5_M13
  `undef AXI_AR_LAYER_S5_M13
`endif 

`ifdef AXI_AR_LAYER_S5_M14
  `undef AXI_AR_LAYER_S5_M14
`endif 

`ifdef AXI_AR_LAYER_S5_M15
  `undef AXI_AR_LAYER_S5_M15
`endif 

`ifdef AXI_AR_LAYER_S5_M16
  `undef AXI_AR_LAYER_S5_M16
`endif 

`ifdef AXI_AW_LAYER_S5_M1
  `undef AXI_AW_LAYER_S5_M1
`endif 

`ifdef AXI_AW_LAYER_S5_M2
  `undef AXI_AW_LAYER_S5_M2
`endif 

`ifdef AXI_AW_LAYER_S5_M3
  `undef AXI_AW_LAYER_S5_M3
`endif 

`ifdef AXI_AW_LAYER_S5_M4
  `undef AXI_AW_LAYER_S5_M4
`endif 

`ifdef AXI_AW_LAYER_S5_M5
  `undef AXI_AW_LAYER_S5_M5
`endif 

`ifdef AXI_AW_LAYER_S5_M6
  `undef AXI_AW_LAYER_S5_M6
`endif 

`ifdef AXI_AW_LAYER_S5_M7
  `undef AXI_AW_LAYER_S5_M7
`endif 

`ifdef AXI_AW_LAYER_S5_M8
  `undef AXI_AW_LAYER_S5_M8
`endif 

`ifdef AXI_AW_LAYER_S5_M9
  `undef AXI_AW_LAYER_S5_M9
`endif 

`ifdef AXI_AW_LAYER_S5_M10
  `undef AXI_AW_LAYER_S5_M10
`endif 

`ifdef AXI_AW_LAYER_S5_M11
  `undef AXI_AW_LAYER_S5_M11
`endif 

`ifdef AXI_AW_LAYER_S5_M12
  `undef AXI_AW_LAYER_S5_M12
`endif 

`ifdef AXI_AW_LAYER_S5_M13
  `undef AXI_AW_LAYER_S5_M13
`endif 

`ifdef AXI_AW_LAYER_S5_M14
  `undef AXI_AW_LAYER_S5_M14
`endif 

`ifdef AXI_AW_LAYER_S5_M15
  `undef AXI_AW_LAYER_S5_M15
`endif 

`ifdef AXI_AW_LAYER_S5_M16
  `undef AXI_AW_LAYER_S5_M16
`endif 

`ifdef AXI_W_LAYER_S5_M1
  `undef AXI_W_LAYER_S5_M1
`endif 

`ifdef AXI_W_LAYER_S5_M2
  `undef AXI_W_LAYER_S5_M2
`endif 

`ifdef AXI_W_LAYER_S5_M3
  `undef AXI_W_LAYER_S5_M3
`endif 

`ifdef AXI_W_LAYER_S5_M4
  `undef AXI_W_LAYER_S5_M4
`endif 

`ifdef AXI_W_LAYER_S5_M5
  `undef AXI_W_LAYER_S5_M5
`endif 

`ifdef AXI_W_LAYER_S5_M6
  `undef AXI_W_LAYER_S5_M6
`endif 

`ifdef AXI_W_LAYER_S5_M7
  `undef AXI_W_LAYER_S5_M7
`endif 

`ifdef AXI_W_LAYER_S5_M8
  `undef AXI_W_LAYER_S5_M8
`endif 

`ifdef AXI_W_LAYER_S5_M9
  `undef AXI_W_LAYER_S5_M9
`endif 

`ifdef AXI_W_LAYER_S5_M10
  `undef AXI_W_LAYER_S5_M10
`endif 

`ifdef AXI_W_LAYER_S5_M11
  `undef AXI_W_LAYER_S5_M11
`endif 

`ifdef AXI_W_LAYER_S5_M12
  `undef AXI_W_LAYER_S5_M12
`endif 

`ifdef AXI_W_LAYER_S5_M13
  `undef AXI_W_LAYER_S5_M13
`endif 

`ifdef AXI_W_LAYER_S5_M14
  `undef AXI_W_LAYER_S5_M14
`endif 

`ifdef AXI_W_LAYER_S5_M15
  `undef AXI_W_LAYER_S5_M15
`endif 

`ifdef AXI_W_LAYER_S5_M16
  `undef AXI_W_LAYER_S5_M16
`endif 

`ifdef AXI_AR_LAYER_S6_M1
  `undef AXI_AR_LAYER_S6_M1
`endif 

`ifdef AXI_AR_LAYER_S6_M2
  `undef AXI_AR_LAYER_S6_M2
`endif 

`ifdef AXI_AR_LAYER_S6_M3
  `undef AXI_AR_LAYER_S6_M3
`endif 

`ifdef AXI_AR_LAYER_S6_M4
  `undef AXI_AR_LAYER_S6_M4
`endif 

`ifdef AXI_AR_LAYER_S6_M5
  `undef AXI_AR_LAYER_S6_M5
`endif 

`ifdef AXI_AR_LAYER_S6_M6
  `undef AXI_AR_LAYER_S6_M6
`endif 

`ifdef AXI_AR_LAYER_S6_M7
  `undef AXI_AR_LAYER_S6_M7
`endif 

`ifdef AXI_AR_LAYER_S6_M8
  `undef AXI_AR_LAYER_S6_M8
`endif 

`ifdef AXI_AR_LAYER_S6_M9
  `undef AXI_AR_LAYER_S6_M9
`endif 

`ifdef AXI_AR_LAYER_S6_M10
  `undef AXI_AR_LAYER_S6_M10
`endif 

`ifdef AXI_AR_LAYER_S6_M11
  `undef AXI_AR_LAYER_S6_M11
`endif 

`ifdef AXI_AR_LAYER_S6_M12
  `undef AXI_AR_LAYER_S6_M12
`endif 

`ifdef AXI_AR_LAYER_S6_M13
  `undef AXI_AR_LAYER_S6_M13
`endif 

`ifdef AXI_AR_LAYER_S6_M14
  `undef AXI_AR_LAYER_S6_M14
`endif 

`ifdef AXI_AR_LAYER_S6_M15
  `undef AXI_AR_LAYER_S6_M15
`endif 

`ifdef AXI_AR_LAYER_S6_M16
  `undef AXI_AR_LAYER_S6_M16
`endif 

`ifdef AXI_AW_LAYER_S6_M1
  `undef AXI_AW_LAYER_S6_M1
`endif 

`ifdef AXI_AW_LAYER_S6_M2
  `undef AXI_AW_LAYER_S6_M2
`endif 

`ifdef AXI_AW_LAYER_S6_M3
  `undef AXI_AW_LAYER_S6_M3
`endif 

`ifdef AXI_AW_LAYER_S6_M4
  `undef AXI_AW_LAYER_S6_M4
`endif 

`ifdef AXI_AW_LAYER_S6_M5
  `undef AXI_AW_LAYER_S6_M5
`endif 

`ifdef AXI_AW_LAYER_S6_M6
  `undef AXI_AW_LAYER_S6_M6
`endif 

`ifdef AXI_AW_LAYER_S6_M7
  `undef AXI_AW_LAYER_S6_M7
`endif 

`ifdef AXI_AW_LAYER_S6_M8
  `undef AXI_AW_LAYER_S6_M8
`endif 

`ifdef AXI_AW_LAYER_S6_M9
  `undef AXI_AW_LAYER_S6_M9
`endif 

`ifdef AXI_AW_LAYER_S6_M10
  `undef AXI_AW_LAYER_S6_M10
`endif 

`ifdef AXI_AW_LAYER_S6_M11
  `undef AXI_AW_LAYER_S6_M11
`endif 

`ifdef AXI_AW_LAYER_S6_M12
  `undef AXI_AW_LAYER_S6_M12
`endif 

`ifdef AXI_AW_LAYER_S6_M13
  `undef AXI_AW_LAYER_S6_M13
`endif 

`ifdef AXI_AW_LAYER_S6_M14
  `undef AXI_AW_LAYER_S6_M14
`endif 

`ifdef AXI_AW_LAYER_S6_M15
  `undef AXI_AW_LAYER_S6_M15
`endif 

`ifdef AXI_AW_LAYER_S6_M16
  `undef AXI_AW_LAYER_S6_M16
`endif 

`ifdef AXI_W_LAYER_S6_M1
  `undef AXI_W_LAYER_S6_M1
`endif 

`ifdef AXI_W_LAYER_S6_M2
  `undef AXI_W_LAYER_S6_M2
`endif 

`ifdef AXI_W_LAYER_S6_M3
  `undef AXI_W_LAYER_S6_M3
`endif 

`ifdef AXI_W_LAYER_S6_M4
  `undef AXI_W_LAYER_S6_M4
`endif 

`ifdef AXI_W_LAYER_S6_M5
  `undef AXI_W_LAYER_S6_M5
`endif 

`ifdef AXI_W_LAYER_S6_M6
  `undef AXI_W_LAYER_S6_M6
`endif 

`ifdef AXI_W_LAYER_S6_M7
  `undef AXI_W_LAYER_S6_M7
`endif 

`ifdef AXI_W_LAYER_S6_M8
  `undef AXI_W_LAYER_S6_M8
`endif 

`ifdef AXI_W_LAYER_S6_M9
  `undef AXI_W_LAYER_S6_M9
`endif 

`ifdef AXI_W_LAYER_S6_M10
  `undef AXI_W_LAYER_S6_M10
`endif 

`ifdef AXI_W_LAYER_S6_M11
  `undef AXI_W_LAYER_S6_M11
`endif 

`ifdef AXI_W_LAYER_S6_M12
  `undef AXI_W_LAYER_S6_M12
`endif 

`ifdef AXI_W_LAYER_S6_M13
  `undef AXI_W_LAYER_S6_M13
`endif 

`ifdef AXI_W_LAYER_S6_M14
  `undef AXI_W_LAYER_S6_M14
`endif 

`ifdef AXI_W_LAYER_S6_M15
  `undef AXI_W_LAYER_S6_M15
`endif 

`ifdef AXI_W_LAYER_S6_M16
  `undef AXI_W_LAYER_S6_M16
`endif 

`ifdef AXI_AR_LAYER_S7_M1
  `undef AXI_AR_LAYER_S7_M1
`endif 

`ifdef AXI_AR_LAYER_S7_M2
  `undef AXI_AR_LAYER_S7_M2
`endif 

`ifdef AXI_AR_LAYER_S7_M3
  `undef AXI_AR_LAYER_S7_M3
`endif 

`ifdef AXI_AR_LAYER_S7_M4
  `undef AXI_AR_LAYER_S7_M4
`endif 

`ifdef AXI_AR_LAYER_S7_M5
  `undef AXI_AR_LAYER_S7_M5
`endif 

`ifdef AXI_AR_LAYER_S7_M6
  `undef AXI_AR_LAYER_S7_M6
`endif 

`ifdef AXI_AR_LAYER_S7_M7
  `undef AXI_AR_LAYER_S7_M7
`endif 

`ifdef AXI_AR_LAYER_S7_M8
  `undef AXI_AR_LAYER_S7_M8
`endif 

`ifdef AXI_AR_LAYER_S7_M9
  `undef AXI_AR_LAYER_S7_M9
`endif 

`ifdef AXI_AR_LAYER_S7_M10
  `undef AXI_AR_LAYER_S7_M10
`endif 

`ifdef AXI_AR_LAYER_S7_M11
  `undef AXI_AR_LAYER_S7_M11
`endif 

`ifdef AXI_AR_LAYER_S7_M12
  `undef AXI_AR_LAYER_S7_M12
`endif 

`ifdef AXI_AR_LAYER_S7_M13
  `undef AXI_AR_LAYER_S7_M13
`endif 

`ifdef AXI_AR_LAYER_S7_M14
  `undef AXI_AR_LAYER_S7_M14
`endif 

`ifdef AXI_AR_LAYER_S7_M15
  `undef AXI_AR_LAYER_S7_M15
`endif 

`ifdef AXI_AR_LAYER_S7_M16
  `undef AXI_AR_LAYER_S7_M16
`endif 

`ifdef AXI_AW_LAYER_S7_M1
  `undef AXI_AW_LAYER_S7_M1
`endif 

`ifdef AXI_AW_LAYER_S7_M2
  `undef AXI_AW_LAYER_S7_M2
`endif 

`ifdef AXI_AW_LAYER_S7_M3
  `undef AXI_AW_LAYER_S7_M3
`endif 

`ifdef AXI_AW_LAYER_S7_M4
  `undef AXI_AW_LAYER_S7_M4
`endif 

`ifdef AXI_AW_LAYER_S7_M5
  `undef AXI_AW_LAYER_S7_M5
`endif 

`ifdef AXI_AW_LAYER_S7_M6
  `undef AXI_AW_LAYER_S7_M6
`endif 

`ifdef AXI_AW_LAYER_S7_M7
  `undef AXI_AW_LAYER_S7_M7
`endif 

`ifdef AXI_AW_LAYER_S7_M8
  `undef AXI_AW_LAYER_S7_M8
`endif 

`ifdef AXI_AW_LAYER_S7_M9
  `undef AXI_AW_LAYER_S7_M9
`endif 

`ifdef AXI_AW_LAYER_S7_M10
  `undef AXI_AW_LAYER_S7_M10
`endif 

`ifdef AXI_AW_LAYER_S7_M11
  `undef AXI_AW_LAYER_S7_M11
`endif 

`ifdef AXI_AW_LAYER_S7_M12
  `undef AXI_AW_LAYER_S7_M12
`endif 

`ifdef AXI_AW_LAYER_S7_M13
  `undef AXI_AW_LAYER_S7_M13
`endif 

`ifdef AXI_AW_LAYER_S7_M14
  `undef AXI_AW_LAYER_S7_M14
`endif 

`ifdef AXI_AW_LAYER_S7_M15
  `undef AXI_AW_LAYER_S7_M15
`endif 

`ifdef AXI_AW_LAYER_S7_M16
  `undef AXI_AW_LAYER_S7_M16
`endif 

`ifdef AXI_W_LAYER_S7_M1
  `undef AXI_W_LAYER_S7_M1
`endif 

`ifdef AXI_W_LAYER_S7_M2
  `undef AXI_W_LAYER_S7_M2
`endif 

`ifdef AXI_W_LAYER_S7_M3
  `undef AXI_W_LAYER_S7_M3
`endif 

`ifdef AXI_W_LAYER_S7_M4
  `undef AXI_W_LAYER_S7_M4
`endif 

`ifdef AXI_W_LAYER_S7_M5
  `undef AXI_W_LAYER_S7_M5
`endif 

`ifdef AXI_W_LAYER_S7_M6
  `undef AXI_W_LAYER_S7_M6
`endif 

`ifdef AXI_W_LAYER_S7_M7
  `undef AXI_W_LAYER_S7_M7
`endif 

`ifdef AXI_W_LAYER_S7_M8
  `undef AXI_W_LAYER_S7_M8
`endif 

`ifdef AXI_W_LAYER_S7_M9
  `undef AXI_W_LAYER_S7_M9
`endif 

`ifdef AXI_W_LAYER_S7_M10
  `undef AXI_W_LAYER_S7_M10
`endif 

`ifdef AXI_W_LAYER_S7_M11
  `undef AXI_W_LAYER_S7_M11
`endif 

`ifdef AXI_W_LAYER_S7_M12
  `undef AXI_W_LAYER_S7_M12
`endif 

`ifdef AXI_W_LAYER_S7_M13
  `undef AXI_W_LAYER_S7_M13
`endif 

`ifdef AXI_W_LAYER_S7_M14
  `undef AXI_W_LAYER_S7_M14
`endif 

`ifdef AXI_W_LAYER_S7_M15
  `undef AXI_W_LAYER_S7_M15
`endif 

`ifdef AXI_W_LAYER_S7_M16
  `undef AXI_W_LAYER_S7_M16
`endif 

`ifdef AXI_AR_LAYER_S8_M1
  `undef AXI_AR_LAYER_S8_M1
`endif 

`ifdef AXI_AR_LAYER_S8_M2
  `undef AXI_AR_LAYER_S8_M2
`endif 

`ifdef AXI_AR_LAYER_S8_M3
  `undef AXI_AR_LAYER_S8_M3
`endif 

`ifdef AXI_AR_LAYER_S8_M4
  `undef AXI_AR_LAYER_S8_M4
`endif 

`ifdef AXI_AR_LAYER_S8_M5
  `undef AXI_AR_LAYER_S8_M5
`endif 

`ifdef AXI_AR_LAYER_S8_M6
  `undef AXI_AR_LAYER_S8_M6
`endif 

`ifdef AXI_AR_LAYER_S8_M7
  `undef AXI_AR_LAYER_S8_M7
`endif 

`ifdef AXI_AR_LAYER_S8_M8
  `undef AXI_AR_LAYER_S8_M8
`endif 

`ifdef AXI_AR_LAYER_S8_M9
  `undef AXI_AR_LAYER_S8_M9
`endif 

`ifdef AXI_AR_LAYER_S8_M10
  `undef AXI_AR_LAYER_S8_M10
`endif 

`ifdef AXI_AR_LAYER_S8_M11
  `undef AXI_AR_LAYER_S8_M11
`endif 

`ifdef AXI_AR_LAYER_S8_M12
  `undef AXI_AR_LAYER_S8_M12
`endif 

`ifdef AXI_AR_LAYER_S8_M13
  `undef AXI_AR_LAYER_S8_M13
`endif 

`ifdef AXI_AR_LAYER_S8_M14
  `undef AXI_AR_LAYER_S8_M14
`endif 

`ifdef AXI_AR_LAYER_S8_M15
  `undef AXI_AR_LAYER_S8_M15
`endif 

`ifdef AXI_AR_LAYER_S8_M16
  `undef AXI_AR_LAYER_S8_M16
`endif 

`ifdef AXI_AW_LAYER_S8_M1
  `undef AXI_AW_LAYER_S8_M1
`endif 

`ifdef AXI_AW_LAYER_S8_M2
  `undef AXI_AW_LAYER_S8_M2
`endif 

`ifdef AXI_AW_LAYER_S8_M3
  `undef AXI_AW_LAYER_S8_M3
`endif 

`ifdef AXI_AW_LAYER_S8_M4
  `undef AXI_AW_LAYER_S8_M4
`endif 

`ifdef AXI_AW_LAYER_S8_M5
  `undef AXI_AW_LAYER_S8_M5
`endif 

`ifdef AXI_AW_LAYER_S8_M6
  `undef AXI_AW_LAYER_S8_M6
`endif 

`ifdef AXI_AW_LAYER_S8_M7
  `undef AXI_AW_LAYER_S8_M7
`endif 

`ifdef AXI_AW_LAYER_S8_M8
  `undef AXI_AW_LAYER_S8_M8
`endif 

`ifdef AXI_AW_LAYER_S8_M9
  `undef AXI_AW_LAYER_S8_M9
`endif 

`ifdef AXI_AW_LAYER_S8_M10
  `undef AXI_AW_LAYER_S8_M10
`endif 

`ifdef AXI_AW_LAYER_S8_M11
  `undef AXI_AW_LAYER_S8_M11
`endif 

`ifdef AXI_AW_LAYER_S8_M12
  `undef AXI_AW_LAYER_S8_M12
`endif 

`ifdef AXI_AW_LAYER_S8_M13
  `undef AXI_AW_LAYER_S8_M13
`endif 

`ifdef AXI_AW_LAYER_S8_M14
  `undef AXI_AW_LAYER_S8_M14
`endif 

`ifdef AXI_AW_LAYER_S8_M15
  `undef AXI_AW_LAYER_S8_M15
`endif 

`ifdef AXI_AW_LAYER_S8_M16
  `undef AXI_AW_LAYER_S8_M16
`endif 

`ifdef AXI_W_LAYER_S8_M1
  `undef AXI_W_LAYER_S8_M1
`endif 

`ifdef AXI_W_LAYER_S8_M2
  `undef AXI_W_LAYER_S8_M2
`endif 

`ifdef AXI_W_LAYER_S8_M3
  `undef AXI_W_LAYER_S8_M3
`endif 

`ifdef AXI_W_LAYER_S8_M4
  `undef AXI_W_LAYER_S8_M4
`endif 

`ifdef AXI_W_LAYER_S8_M5
  `undef AXI_W_LAYER_S8_M5
`endif 

`ifdef AXI_W_LAYER_S8_M6
  `undef AXI_W_LAYER_S8_M6
`endif 

`ifdef AXI_W_LAYER_S8_M7
  `undef AXI_W_LAYER_S8_M7
`endif 

`ifdef AXI_W_LAYER_S8_M8
  `undef AXI_W_LAYER_S8_M8
`endif 

`ifdef AXI_W_LAYER_S8_M9
  `undef AXI_W_LAYER_S8_M9
`endif 

`ifdef AXI_W_LAYER_S8_M10
  `undef AXI_W_LAYER_S8_M10
`endif 

`ifdef AXI_W_LAYER_S8_M11
  `undef AXI_W_LAYER_S8_M11
`endif 

`ifdef AXI_W_LAYER_S8_M12
  `undef AXI_W_LAYER_S8_M12
`endif 

`ifdef AXI_W_LAYER_S8_M13
  `undef AXI_W_LAYER_S8_M13
`endif 

`ifdef AXI_W_LAYER_S8_M14
  `undef AXI_W_LAYER_S8_M14
`endif 

`ifdef AXI_W_LAYER_S8_M15
  `undef AXI_W_LAYER_S8_M15
`endif 

`ifdef AXI_W_LAYER_S8_M16
  `undef AXI_W_LAYER_S8_M16
`endif 

`ifdef AXI_AR_LAYER_S9_M1
  `undef AXI_AR_LAYER_S9_M1
`endif 

`ifdef AXI_AR_LAYER_S9_M2
  `undef AXI_AR_LAYER_S9_M2
`endif 

`ifdef AXI_AR_LAYER_S9_M3
  `undef AXI_AR_LAYER_S9_M3
`endif 

`ifdef AXI_AR_LAYER_S9_M4
  `undef AXI_AR_LAYER_S9_M4
`endif 

`ifdef AXI_AR_LAYER_S9_M5
  `undef AXI_AR_LAYER_S9_M5
`endif 

`ifdef AXI_AR_LAYER_S9_M6
  `undef AXI_AR_LAYER_S9_M6
`endif 

`ifdef AXI_AR_LAYER_S9_M7
  `undef AXI_AR_LAYER_S9_M7
`endif 

`ifdef AXI_AR_LAYER_S9_M8
  `undef AXI_AR_LAYER_S9_M8
`endif 

`ifdef AXI_AR_LAYER_S9_M9
  `undef AXI_AR_LAYER_S9_M9
`endif 

`ifdef AXI_AR_LAYER_S9_M10
  `undef AXI_AR_LAYER_S9_M10
`endif 

`ifdef AXI_AR_LAYER_S9_M11
  `undef AXI_AR_LAYER_S9_M11
`endif 

`ifdef AXI_AR_LAYER_S9_M12
  `undef AXI_AR_LAYER_S9_M12
`endif 

`ifdef AXI_AR_LAYER_S9_M13
  `undef AXI_AR_LAYER_S9_M13
`endif 

`ifdef AXI_AR_LAYER_S9_M14
  `undef AXI_AR_LAYER_S9_M14
`endif 

`ifdef AXI_AR_LAYER_S9_M15
  `undef AXI_AR_LAYER_S9_M15
`endif 

`ifdef AXI_AR_LAYER_S9_M16
  `undef AXI_AR_LAYER_S9_M16
`endif 

`ifdef AXI_AW_LAYER_S9_M1
  `undef AXI_AW_LAYER_S9_M1
`endif 

`ifdef AXI_AW_LAYER_S9_M2
  `undef AXI_AW_LAYER_S9_M2
`endif 

`ifdef AXI_AW_LAYER_S9_M3
  `undef AXI_AW_LAYER_S9_M3
`endif 

`ifdef AXI_AW_LAYER_S9_M4
  `undef AXI_AW_LAYER_S9_M4
`endif 

`ifdef AXI_AW_LAYER_S9_M5
  `undef AXI_AW_LAYER_S9_M5
`endif 

`ifdef AXI_AW_LAYER_S9_M6
  `undef AXI_AW_LAYER_S9_M6
`endif 

`ifdef AXI_AW_LAYER_S9_M7
  `undef AXI_AW_LAYER_S9_M7
`endif 

`ifdef AXI_AW_LAYER_S9_M8
  `undef AXI_AW_LAYER_S9_M8
`endif 

`ifdef AXI_AW_LAYER_S9_M9
  `undef AXI_AW_LAYER_S9_M9
`endif 

`ifdef AXI_AW_LAYER_S9_M10
  `undef AXI_AW_LAYER_S9_M10
`endif 

`ifdef AXI_AW_LAYER_S9_M11
  `undef AXI_AW_LAYER_S9_M11
`endif 

`ifdef AXI_AW_LAYER_S9_M12
  `undef AXI_AW_LAYER_S9_M12
`endif 

`ifdef AXI_AW_LAYER_S9_M13
  `undef AXI_AW_LAYER_S9_M13
`endif 

`ifdef AXI_AW_LAYER_S9_M14
  `undef AXI_AW_LAYER_S9_M14
`endif 

`ifdef AXI_AW_LAYER_S9_M15
  `undef AXI_AW_LAYER_S9_M15
`endif 

`ifdef AXI_AW_LAYER_S9_M16
  `undef AXI_AW_LAYER_S9_M16
`endif 

`ifdef AXI_W_LAYER_S9_M1
  `undef AXI_W_LAYER_S9_M1
`endif 

`ifdef AXI_W_LAYER_S9_M2
  `undef AXI_W_LAYER_S9_M2
`endif 

`ifdef AXI_W_LAYER_S9_M3
  `undef AXI_W_LAYER_S9_M3
`endif 

`ifdef AXI_W_LAYER_S9_M4
  `undef AXI_W_LAYER_S9_M4
`endif 

`ifdef AXI_W_LAYER_S9_M5
  `undef AXI_W_LAYER_S9_M5
`endif 

`ifdef AXI_W_LAYER_S9_M6
  `undef AXI_W_LAYER_S9_M6
`endif 

`ifdef AXI_W_LAYER_S9_M7
  `undef AXI_W_LAYER_S9_M7
`endif 

`ifdef AXI_W_LAYER_S9_M8
  `undef AXI_W_LAYER_S9_M8
`endif 

`ifdef AXI_W_LAYER_S9_M9
  `undef AXI_W_LAYER_S9_M9
`endif 

`ifdef AXI_W_LAYER_S9_M10
  `undef AXI_W_LAYER_S9_M10
`endif 

`ifdef AXI_W_LAYER_S9_M11
  `undef AXI_W_LAYER_S9_M11
`endif 

`ifdef AXI_W_LAYER_S9_M12
  `undef AXI_W_LAYER_S9_M12
`endif 

`ifdef AXI_W_LAYER_S9_M13
  `undef AXI_W_LAYER_S9_M13
`endif 

`ifdef AXI_W_LAYER_S9_M14
  `undef AXI_W_LAYER_S9_M14
`endif 

`ifdef AXI_W_LAYER_S9_M15
  `undef AXI_W_LAYER_S9_M15
`endif 

`ifdef AXI_W_LAYER_S9_M16
  `undef AXI_W_LAYER_S9_M16
`endif 

`ifdef AXI_AR_LAYER_S10_M1
  `undef AXI_AR_LAYER_S10_M1
`endif 

`ifdef AXI_AR_LAYER_S10_M2
  `undef AXI_AR_LAYER_S10_M2
`endif 

`ifdef AXI_AR_LAYER_S10_M3
  `undef AXI_AR_LAYER_S10_M3
`endif 

`ifdef AXI_AR_LAYER_S10_M4
  `undef AXI_AR_LAYER_S10_M4
`endif 

`ifdef AXI_AR_LAYER_S10_M5
  `undef AXI_AR_LAYER_S10_M5
`endif 

`ifdef AXI_AR_LAYER_S10_M6
  `undef AXI_AR_LAYER_S10_M6
`endif 

`ifdef AXI_AR_LAYER_S10_M7
  `undef AXI_AR_LAYER_S10_M7
`endif 

`ifdef AXI_AR_LAYER_S10_M8
  `undef AXI_AR_LAYER_S10_M8
`endif 

`ifdef AXI_AR_LAYER_S10_M9
  `undef AXI_AR_LAYER_S10_M9
`endif 

`ifdef AXI_AR_LAYER_S10_M10
  `undef AXI_AR_LAYER_S10_M10
`endif 

`ifdef AXI_AR_LAYER_S10_M11
  `undef AXI_AR_LAYER_S10_M11
`endif 

`ifdef AXI_AR_LAYER_S10_M12
  `undef AXI_AR_LAYER_S10_M12
`endif 

`ifdef AXI_AR_LAYER_S10_M13
  `undef AXI_AR_LAYER_S10_M13
`endif 

`ifdef AXI_AR_LAYER_S10_M14
  `undef AXI_AR_LAYER_S10_M14
`endif 

`ifdef AXI_AR_LAYER_S10_M15
  `undef AXI_AR_LAYER_S10_M15
`endif 

`ifdef AXI_AR_LAYER_S10_M16
  `undef AXI_AR_LAYER_S10_M16
`endif 

`ifdef AXI_AW_LAYER_S10_M1
  `undef AXI_AW_LAYER_S10_M1
`endif 

`ifdef AXI_AW_LAYER_S10_M2
  `undef AXI_AW_LAYER_S10_M2
`endif 

`ifdef AXI_AW_LAYER_S10_M3
  `undef AXI_AW_LAYER_S10_M3
`endif 

`ifdef AXI_AW_LAYER_S10_M4
  `undef AXI_AW_LAYER_S10_M4
`endif 

`ifdef AXI_AW_LAYER_S10_M5
  `undef AXI_AW_LAYER_S10_M5
`endif 

`ifdef AXI_AW_LAYER_S10_M6
  `undef AXI_AW_LAYER_S10_M6
`endif 

`ifdef AXI_AW_LAYER_S10_M7
  `undef AXI_AW_LAYER_S10_M7
`endif 

`ifdef AXI_AW_LAYER_S10_M8
  `undef AXI_AW_LAYER_S10_M8
`endif 

`ifdef AXI_AW_LAYER_S10_M9
  `undef AXI_AW_LAYER_S10_M9
`endif 

`ifdef AXI_AW_LAYER_S10_M10
  `undef AXI_AW_LAYER_S10_M10
`endif 

`ifdef AXI_AW_LAYER_S10_M11
  `undef AXI_AW_LAYER_S10_M11
`endif 

`ifdef AXI_AW_LAYER_S10_M12
  `undef AXI_AW_LAYER_S10_M12
`endif 

`ifdef AXI_AW_LAYER_S10_M13
  `undef AXI_AW_LAYER_S10_M13
`endif 

`ifdef AXI_AW_LAYER_S10_M14
  `undef AXI_AW_LAYER_S10_M14
`endif 

`ifdef AXI_AW_LAYER_S10_M15
  `undef AXI_AW_LAYER_S10_M15
`endif 

`ifdef AXI_AW_LAYER_S10_M16
  `undef AXI_AW_LAYER_S10_M16
`endif 

`ifdef AXI_W_LAYER_S10_M1
  `undef AXI_W_LAYER_S10_M1
`endif 

`ifdef AXI_W_LAYER_S10_M2
  `undef AXI_W_LAYER_S10_M2
`endif 

`ifdef AXI_W_LAYER_S10_M3
  `undef AXI_W_LAYER_S10_M3
`endif 

`ifdef AXI_W_LAYER_S10_M4
  `undef AXI_W_LAYER_S10_M4
`endif 

`ifdef AXI_W_LAYER_S10_M5
  `undef AXI_W_LAYER_S10_M5
`endif 

`ifdef AXI_W_LAYER_S10_M6
  `undef AXI_W_LAYER_S10_M6
`endif 

`ifdef AXI_W_LAYER_S10_M7
  `undef AXI_W_LAYER_S10_M7
`endif 

`ifdef AXI_W_LAYER_S10_M8
  `undef AXI_W_LAYER_S10_M8
`endif 

`ifdef AXI_W_LAYER_S10_M9
  `undef AXI_W_LAYER_S10_M9
`endif 

`ifdef AXI_W_LAYER_S10_M10
  `undef AXI_W_LAYER_S10_M10
`endif 

`ifdef AXI_W_LAYER_S10_M11
  `undef AXI_W_LAYER_S10_M11
`endif 

`ifdef AXI_W_LAYER_S10_M12
  `undef AXI_W_LAYER_S10_M12
`endif 

`ifdef AXI_W_LAYER_S10_M13
  `undef AXI_W_LAYER_S10_M13
`endif 

`ifdef AXI_W_LAYER_S10_M14
  `undef AXI_W_LAYER_S10_M14
`endif 

`ifdef AXI_W_LAYER_S10_M15
  `undef AXI_W_LAYER_S10_M15
`endif 

`ifdef AXI_W_LAYER_S10_M16
  `undef AXI_W_LAYER_S10_M16
`endif 

`ifdef AXI_AR_LAYER_S11_M1
  `undef AXI_AR_LAYER_S11_M1
`endif 

`ifdef AXI_AR_LAYER_S11_M2
  `undef AXI_AR_LAYER_S11_M2
`endif 

`ifdef AXI_AR_LAYER_S11_M3
  `undef AXI_AR_LAYER_S11_M3
`endif 

`ifdef AXI_AR_LAYER_S11_M4
  `undef AXI_AR_LAYER_S11_M4
`endif 

`ifdef AXI_AR_LAYER_S11_M5
  `undef AXI_AR_LAYER_S11_M5
`endif 

`ifdef AXI_AR_LAYER_S11_M6
  `undef AXI_AR_LAYER_S11_M6
`endif 

`ifdef AXI_AR_LAYER_S11_M7
  `undef AXI_AR_LAYER_S11_M7
`endif 

`ifdef AXI_AR_LAYER_S11_M8
  `undef AXI_AR_LAYER_S11_M8
`endif 

`ifdef AXI_AR_LAYER_S11_M9
  `undef AXI_AR_LAYER_S11_M9
`endif 

`ifdef AXI_AR_LAYER_S11_M10
  `undef AXI_AR_LAYER_S11_M10
`endif 

`ifdef AXI_AR_LAYER_S11_M11
  `undef AXI_AR_LAYER_S11_M11
`endif 

`ifdef AXI_AR_LAYER_S11_M12
  `undef AXI_AR_LAYER_S11_M12
`endif 

`ifdef AXI_AR_LAYER_S11_M13
  `undef AXI_AR_LAYER_S11_M13
`endif 

`ifdef AXI_AR_LAYER_S11_M14
  `undef AXI_AR_LAYER_S11_M14
`endif 

`ifdef AXI_AR_LAYER_S11_M15
  `undef AXI_AR_LAYER_S11_M15
`endif 

`ifdef AXI_AR_LAYER_S11_M16
  `undef AXI_AR_LAYER_S11_M16
`endif 

`ifdef AXI_AW_LAYER_S11_M1
  `undef AXI_AW_LAYER_S11_M1
`endif 

`ifdef AXI_AW_LAYER_S11_M2
  `undef AXI_AW_LAYER_S11_M2
`endif 

`ifdef AXI_AW_LAYER_S11_M3
  `undef AXI_AW_LAYER_S11_M3
`endif 

`ifdef AXI_AW_LAYER_S11_M4
  `undef AXI_AW_LAYER_S11_M4
`endif 

`ifdef AXI_AW_LAYER_S11_M5
  `undef AXI_AW_LAYER_S11_M5
`endif 

`ifdef AXI_AW_LAYER_S11_M6
  `undef AXI_AW_LAYER_S11_M6
`endif 

`ifdef AXI_AW_LAYER_S11_M7
  `undef AXI_AW_LAYER_S11_M7
`endif 

`ifdef AXI_AW_LAYER_S11_M8
  `undef AXI_AW_LAYER_S11_M8
`endif 

`ifdef AXI_AW_LAYER_S11_M9
  `undef AXI_AW_LAYER_S11_M9
`endif 

`ifdef AXI_AW_LAYER_S11_M10
  `undef AXI_AW_LAYER_S11_M10
`endif 

`ifdef AXI_AW_LAYER_S11_M11
  `undef AXI_AW_LAYER_S11_M11
`endif 

`ifdef AXI_AW_LAYER_S11_M12
  `undef AXI_AW_LAYER_S11_M12
`endif 

`ifdef AXI_AW_LAYER_S11_M13
  `undef AXI_AW_LAYER_S11_M13
`endif 

`ifdef AXI_AW_LAYER_S11_M14
  `undef AXI_AW_LAYER_S11_M14
`endif 

`ifdef AXI_AW_LAYER_S11_M15
  `undef AXI_AW_LAYER_S11_M15
`endif 

`ifdef AXI_AW_LAYER_S11_M16
  `undef AXI_AW_LAYER_S11_M16
`endif 

`ifdef AXI_W_LAYER_S11_M1
  `undef AXI_W_LAYER_S11_M1
`endif 

`ifdef AXI_W_LAYER_S11_M2
  `undef AXI_W_LAYER_S11_M2
`endif 

`ifdef AXI_W_LAYER_S11_M3
  `undef AXI_W_LAYER_S11_M3
`endif 

`ifdef AXI_W_LAYER_S11_M4
  `undef AXI_W_LAYER_S11_M4
`endif 

`ifdef AXI_W_LAYER_S11_M5
  `undef AXI_W_LAYER_S11_M5
`endif 

`ifdef AXI_W_LAYER_S11_M6
  `undef AXI_W_LAYER_S11_M6
`endif 

`ifdef AXI_W_LAYER_S11_M7
  `undef AXI_W_LAYER_S11_M7
`endif 

`ifdef AXI_W_LAYER_S11_M8
  `undef AXI_W_LAYER_S11_M8
`endif 

`ifdef AXI_W_LAYER_S11_M9
  `undef AXI_W_LAYER_S11_M9
`endif 

`ifdef AXI_W_LAYER_S11_M10
  `undef AXI_W_LAYER_S11_M10
`endif 

`ifdef AXI_W_LAYER_S11_M11
  `undef AXI_W_LAYER_S11_M11
`endif 

`ifdef AXI_W_LAYER_S11_M12
  `undef AXI_W_LAYER_S11_M12
`endif 

`ifdef AXI_W_LAYER_S11_M13
  `undef AXI_W_LAYER_S11_M13
`endif 

`ifdef AXI_W_LAYER_S11_M14
  `undef AXI_W_LAYER_S11_M14
`endif 

`ifdef AXI_W_LAYER_S11_M15
  `undef AXI_W_LAYER_S11_M15
`endif 

`ifdef AXI_W_LAYER_S11_M16
  `undef AXI_W_LAYER_S11_M16
`endif 

`ifdef AXI_AR_LAYER_S12_M1
  `undef AXI_AR_LAYER_S12_M1
`endif 

`ifdef AXI_AR_LAYER_S12_M2
  `undef AXI_AR_LAYER_S12_M2
`endif 

`ifdef AXI_AR_LAYER_S12_M3
  `undef AXI_AR_LAYER_S12_M3
`endif 

`ifdef AXI_AR_LAYER_S12_M4
  `undef AXI_AR_LAYER_S12_M4
`endif 

`ifdef AXI_AR_LAYER_S12_M5
  `undef AXI_AR_LAYER_S12_M5
`endif 

`ifdef AXI_AR_LAYER_S12_M6
  `undef AXI_AR_LAYER_S12_M6
`endif 

`ifdef AXI_AR_LAYER_S12_M7
  `undef AXI_AR_LAYER_S12_M7
`endif 

`ifdef AXI_AR_LAYER_S12_M8
  `undef AXI_AR_LAYER_S12_M8
`endif 

`ifdef AXI_AR_LAYER_S12_M9
  `undef AXI_AR_LAYER_S12_M9
`endif 

`ifdef AXI_AR_LAYER_S12_M10
  `undef AXI_AR_LAYER_S12_M10
`endif 

`ifdef AXI_AR_LAYER_S12_M11
  `undef AXI_AR_LAYER_S12_M11
`endif 

`ifdef AXI_AR_LAYER_S12_M12
  `undef AXI_AR_LAYER_S12_M12
`endif 

`ifdef AXI_AR_LAYER_S12_M13
  `undef AXI_AR_LAYER_S12_M13
`endif 

`ifdef AXI_AR_LAYER_S12_M14
  `undef AXI_AR_LAYER_S12_M14
`endif 

`ifdef AXI_AR_LAYER_S12_M15
  `undef AXI_AR_LAYER_S12_M15
`endif 

`ifdef AXI_AR_LAYER_S12_M16
  `undef AXI_AR_LAYER_S12_M16
`endif 

`ifdef AXI_AW_LAYER_S12_M1
  `undef AXI_AW_LAYER_S12_M1
`endif 

`ifdef AXI_AW_LAYER_S12_M2
  `undef AXI_AW_LAYER_S12_M2
`endif 

`ifdef AXI_AW_LAYER_S12_M3
  `undef AXI_AW_LAYER_S12_M3
`endif 

`ifdef AXI_AW_LAYER_S12_M4
  `undef AXI_AW_LAYER_S12_M4
`endif 

`ifdef AXI_AW_LAYER_S12_M5
  `undef AXI_AW_LAYER_S12_M5
`endif 

`ifdef AXI_AW_LAYER_S12_M6
  `undef AXI_AW_LAYER_S12_M6
`endif 

`ifdef AXI_AW_LAYER_S12_M7
  `undef AXI_AW_LAYER_S12_M7
`endif 

`ifdef AXI_AW_LAYER_S12_M8
  `undef AXI_AW_LAYER_S12_M8
`endif 

`ifdef AXI_AW_LAYER_S12_M9
  `undef AXI_AW_LAYER_S12_M9
`endif 

`ifdef AXI_AW_LAYER_S12_M10
  `undef AXI_AW_LAYER_S12_M10
`endif 

`ifdef AXI_AW_LAYER_S12_M11
  `undef AXI_AW_LAYER_S12_M11
`endif 

`ifdef AXI_AW_LAYER_S12_M12
  `undef AXI_AW_LAYER_S12_M12
`endif 

`ifdef AXI_AW_LAYER_S12_M13
  `undef AXI_AW_LAYER_S12_M13
`endif 

`ifdef AXI_AW_LAYER_S12_M14
  `undef AXI_AW_LAYER_S12_M14
`endif 

`ifdef AXI_AW_LAYER_S12_M15
  `undef AXI_AW_LAYER_S12_M15
`endif 

`ifdef AXI_AW_LAYER_S12_M16
  `undef AXI_AW_LAYER_S12_M16
`endif 

`ifdef AXI_W_LAYER_S12_M1
  `undef AXI_W_LAYER_S12_M1
`endif 

`ifdef AXI_W_LAYER_S12_M2
  `undef AXI_W_LAYER_S12_M2
`endif 

`ifdef AXI_W_LAYER_S12_M3
  `undef AXI_W_LAYER_S12_M3
`endif 

`ifdef AXI_W_LAYER_S12_M4
  `undef AXI_W_LAYER_S12_M4
`endif 

`ifdef AXI_W_LAYER_S12_M5
  `undef AXI_W_LAYER_S12_M5
`endif 

`ifdef AXI_W_LAYER_S12_M6
  `undef AXI_W_LAYER_S12_M6
`endif 

`ifdef AXI_W_LAYER_S12_M7
  `undef AXI_W_LAYER_S12_M7
`endif 

`ifdef AXI_W_LAYER_S12_M8
  `undef AXI_W_LAYER_S12_M8
`endif 

`ifdef AXI_W_LAYER_S12_M9
  `undef AXI_W_LAYER_S12_M9
`endif 

`ifdef AXI_W_LAYER_S12_M10
  `undef AXI_W_LAYER_S12_M10
`endif 

`ifdef AXI_W_LAYER_S12_M11
  `undef AXI_W_LAYER_S12_M11
`endif 

`ifdef AXI_W_LAYER_S12_M12
  `undef AXI_W_LAYER_S12_M12
`endif 

`ifdef AXI_W_LAYER_S12_M13
  `undef AXI_W_LAYER_S12_M13
`endif 

`ifdef AXI_W_LAYER_S12_M14
  `undef AXI_W_LAYER_S12_M14
`endif 

`ifdef AXI_W_LAYER_S12_M15
  `undef AXI_W_LAYER_S12_M15
`endif 

`ifdef AXI_W_LAYER_S12_M16
  `undef AXI_W_LAYER_S12_M16
`endif 

`ifdef AXI_AR_LAYER_S13_M1
  `undef AXI_AR_LAYER_S13_M1
`endif 

`ifdef AXI_AR_LAYER_S13_M2
  `undef AXI_AR_LAYER_S13_M2
`endif 

`ifdef AXI_AR_LAYER_S13_M3
  `undef AXI_AR_LAYER_S13_M3
`endif 

`ifdef AXI_AR_LAYER_S13_M4
  `undef AXI_AR_LAYER_S13_M4
`endif 

`ifdef AXI_AR_LAYER_S13_M5
  `undef AXI_AR_LAYER_S13_M5
`endif 

`ifdef AXI_AR_LAYER_S13_M6
  `undef AXI_AR_LAYER_S13_M6
`endif 

`ifdef AXI_AR_LAYER_S13_M7
  `undef AXI_AR_LAYER_S13_M7
`endif 

`ifdef AXI_AR_LAYER_S13_M8
  `undef AXI_AR_LAYER_S13_M8
`endif 

`ifdef AXI_AR_LAYER_S13_M9
  `undef AXI_AR_LAYER_S13_M9
`endif 

`ifdef AXI_AR_LAYER_S13_M10
  `undef AXI_AR_LAYER_S13_M10
`endif 

`ifdef AXI_AR_LAYER_S13_M11
  `undef AXI_AR_LAYER_S13_M11
`endif 

`ifdef AXI_AR_LAYER_S13_M12
  `undef AXI_AR_LAYER_S13_M12
`endif 

`ifdef AXI_AR_LAYER_S13_M13
  `undef AXI_AR_LAYER_S13_M13
`endif 

`ifdef AXI_AR_LAYER_S13_M14
  `undef AXI_AR_LAYER_S13_M14
`endif 

`ifdef AXI_AR_LAYER_S13_M15
  `undef AXI_AR_LAYER_S13_M15
`endif 

`ifdef AXI_AR_LAYER_S13_M16
  `undef AXI_AR_LAYER_S13_M16
`endif 

`ifdef AXI_AW_LAYER_S13_M1
  `undef AXI_AW_LAYER_S13_M1
`endif 

`ifdef AXI_AW_LAYER_S13_M2
  `undef AXI_AW_LAYER_S13_M2
`endif 

`ifdef AXI_AW_LAYER_S13_M3
  `undef AXI_AW_LAYER_S13_M3
`endif 

`ifdef AXI_AW_LAYER_S13_M4
  `undef AXI_AW_LAYER_S13_M4
`endif 

`ifdef AXI_AW_LAYER_S13_M5
  `undef AXI_AW_LAYER_S13_M5
`endif 

`ifdef AXI_AW_LAYER_S13_M6
  `undef AXI_AW_LAYER_S13_M6
`endif 

`ifdef AXI_AW_LAYER_S13_M7
  `undef AXI_AW_LAYER_S13_M7
`endif 

`ifdef AXI_AW_LAYER_S13_M8
  `undef AXI_AW_LAYER_S13_M8
`endif 

`ifdef AXI_AW_LAYER_S13_M9
  `undef AXI_AW_LAYER_S13_M9
`endif 

`ifdef AXI_AW_LAYER_S13_M10
  `undef AXI_AW_LAYER_S13_M10
`endif 

`ifdef AXI_AW_LAYER_S13_M11
  `undef AXI_AW_LAYER_S13_M11
`endif 

`ifdef AXI_AW_LAYER_S13_M12
  `undef AXI_AW_LAYER_S13_M12
`endif 

`ifdef AXI_AW_LAYER_S13_M13
  `undef AXI_AW_LAYER_S13_M13
`endif 

`ifdef AXI_AW_LAYER_S13_M14
  `undef AXI_AW_LAYER_S13_M14
`endif 

`ifdef AXI_AW_LAYER_S13_M15
  `undef AXI_AW_LAYER_S13_M15
`endif 

`ifdef AXI_AW_LAYER_S13_M16
  `undef AXI_AW_LAYER_S13_M16
`endif 

`ifdef AXI_W_LAYER_S13_M1
  `undef AXI_W_LAYER_S13_M1
`endif 

`ifdef AXI_W_LAYER_S13_M2
  `undef AXI_W_LAYER_S13_M2
`endif 

`ifdef AXI_W_LAYER_S13_M3
  `undef AXI_W_LAYER_S13_M3
`endif 

`ifdef AXI_W_LAYER_S13_M4
  `undef AXI_W_LAYER_S13_M4
`endif 

`ifdef AXI_W_LAYER_S13_M5
  `undef AXI_W_LAYER_S13_M5
`endif 

`ifdef AXI_W_LAYER_S13_M6
  `undef AXI_W_LAYER_S13_M6
`endif 

`ifdef AXI_W_LAYER_S13_M7
  `undef AXI_W_LAYER_S13_M7
`endif 

`ifdef AXI_W_LAYER_S13_M8
  `undef AXI_W_LAYER_S13_M8
`endif 

`ifdef AXI_W_LAYER_S13_M9
  `undef AXI_W_LAYER_S13_M9
`endif 

`ifdef AXI_W_LAYER_S13_M10
  `undef AXI_W_LAYER_S13_M10
`endif 

`ifdef AXI_W_LAYER_S13_M11
  `undef AXI_W_LAYER_S13_M11
`endif 

`ifdef AXI_W_LAYER_S13_M12
  `undef AXI_W_LAYER_S13_M12
`endif 

`ifdef AXI_W_LAYER_S13_M13
  `undef AXI_W_LAYER_S13_M13
`endif 

`ifdef AXI_W_LAYER_S13_M14
  `undef AXI_W_LAYER_S13_M14
`endif 

`ifdef AXI_W_LAYER_S13_M15
  `undef AXI_W_LAYER_S13_M15
`endif 

`ifdef AXI_W_LAYER_S13_M16
  `undef AXI_W_LAYER_S13_M16
`endif 

`ifdef AXI_AR_LAYER_S14_M1
  `undef AXI_AR_LAYER_S14_M1
`endif 

`ifdef AXI_AR_LAYER_S14_M2
  `undef AXI_AR_LAYER_S14_M2
`endif 

`ifdef AXI_AR_LAYER_S14_M3
  `undef AXI_AR_LAYER_S14_M3
`endif 

`ifdef AXI_AR_LAYER_S14_M4
  `undef AXI_AR_LAYER_S14_M4
`endif 

`ifdef AXI_AR_LAYER_S14_M5
  `undef AXI_AR_LAYER_S14_M5
`endif 

`ifdef AXI_AR_LAYER_S14_M6
  `undef AXI_AR_LAYER_S14_M6
`endif 

`ifdef AXI_AR_LAYER_S14_M7
  `undef AXI_AR_LAYER_S14_M7
`endif 

`ifdef AXI_AR_LAYER_S14_M8
  `undef AXI_AR_LAYER_S14_M8
`endif 

`ifdef AXI_AR_LAYER_S14_M9
  `undef AXI_AR_LAYER_S14_M9
`endif 

`ifdef AXI_AR_LAYER_S14_M10
  `undef AXI_AR_LAYER_S14_M10
`endif 

`ifdef AXI_AR_LAYER_S14_M11
  `undef AXI_AR_LAYER_S14_M11
`endif 

`ifdef AXI_AR_LAYER_S14_M12
  `undef AXI_AR_LAYER_S14_M12
`endif 

`ifdef AXI_AR_LAYER_S14_M13
  `undef AXI_AR_LAYER_S14_M13
`endif 

`ifdef AXI_AR_LAYER_S14_M14
  `undef AXI_AR_LAYER_S14_M14
`endif 

`ifdef AXI_AR_LAYER_S14_M15
  `undef AXI_AR_LAYER_S14_M15
`endif 

`ifdef AXI_AR_LAYER_S14_M16
  `undef AXI_AR_LAYER_S14_M16
`endif 

`ifdef AXI_AW_LAYER_S14_M1
  `undef AXI_AW_LAYER_S14_M1
`endif 

`ifdef AXI_AW_LAYER_S14_M2
  `undef AXI_AW_LAYER_S14_M2
`endif 

`ifdef AXI_AW_LAYER_S14_M3
  `undef AXI_AW_LAYER_S14_M3
`endif 

`ifdef AXI_AW_LAYER_S14_M4
  `undef AXI_AW_LAYER_S14_M4
`endif 

`ifdef AXI_AW_LAYER_S14_M5
  `undef AXI_AW_LAYER_S14_M5
`endif 

`ifdef AXI_AW_LAYER_S14_M6
  `undef AXI_AW_LAYER_S14_M6
`endif 

`ifdef AXI_AW_LAYER_S14_M7
  `undef AXI_AW_LAYER_S14_M7
`endif 

`ifdef AXI_AW_LAYER_S14_M8
  `undef AXI_AW_LAYER_S14_M8
`endif 

`ifdef AXI_AW_LAYER_S14_M9
  `undef AXI_AW_LAYER_S14_M9
`endif 

`ifdef AXI_AW_LAYER_S14_M10
  `undef AXI_AW_LAYER_S14_M10
`endif 

`ifdef AXI_AW_LAYER_S14_M11
  `undef AXI_AW_LAYER_S14_M11
`endif 

`ifdef AXI_AW_LAYER_S14_M12
  `undef AXI_AW_LAYER_S14_M12
`endif 

`ifdef AXI_AW_LAYER_S14_M13
  `undef AXI_AW_LAYER_S14_M13
`endif 

`ifdef AXI_AW_LAYER_S14_M14
  `undef AXI_AW_LAYER_S14_M14
`endif 

`ifdef AXI_AW_LAYER_S14_M15
  `undef AXI_AW_LAYER_S14_M15
`endif 

`ifdef AXI_AW_LAYER_S14_M16
  `undef AXI_AW_LAYER_S14_M16
`endif 

`ifdef AXI_W_LAYER_S14_M1
  `undef AXI_W_LAYER_S14_M1
`endif 

`ifdef AXI_W_LAYER_S14_M2
  `undef AXI_W_LAYER_S14_M2
`endif 

`ifdef AXI_W_LAYER_S14_M3
  `undef AXI_W_LAYER_S14_M3
`endif 

`ifdef AXI_W_LAYER_S14_M4
  `undef AXI_W_LAYER_S14_M4
`endif 

`ifdef AXI_W_LAYER_S14_M5
  `undef AXI_W_LAYER_S14_M5
`endif 

`ifdef AXI_W_LAYER_S14_M6
  `undef AXI_W_LAYER_S14_M6
`endif 

`ifdef AXI_W_LAYER_S14_M7
  `undef AXI_W_LAYER_S14_M7
`endif 

`ifdef AXI_W_LAYER_S14_M8
  `undef AXI_W_LAYER_S14_M8
`endif 

`ifdef AXI_W_LAYER_S14_M9
  `undef AXI_W_LAYER_S14_M9
`endif 

`ifdef AXI_W_LAYER_S14_M10
  `undef AXI_W_LAYER_S14_M10
`endif 

`ifdef AXI_W_LAYER_S14_M11
  `undef AXI_W_LAYER_S14_M11
`endif 

`ifdef AXI_W_LAYER_S14_M12
  `undef AXI_W_LAYER_S14_M12
`endif 

`ifdef AXI_W_LAYER_S14_M13
  `undef AXI_W_LAYER_S14_M13
`endif 

`ifdef AXI_W_LAYER_S14_M14
  `undef AXI_W_LAYER_S14_M14
`endif 

`ifdef AXI_W_LAYER_S14_M15
  `undef AXI_W_LAYER_S14_M15
`endif 

`ifdef AXI_W_LAYER_S14_M16
  `undef AXI_W_LAYER_S14_M16
`endif 

`ifdef AXI_AR_LAYER_S15_M1
  `undef AXI_AR_LAYER_S15_M1
`endif 

`ifdef AXI_AR_LAYER_S15_M2
  `undef AXI_AR_LAYER_S15_M2
`endif 

`ifdef AXI_AR_LAYER_S15_M3
  `undef AXI_AR_LAYER_S15_M3
`endif 

`ifdef AXI_AR_LAYER_S15_M4
  `undef AXI_AR_LAYER_S15_M4
`endif 

`ifdef AXI_AR_LAYER_S15_M5
  `undef AXI_AR_LAYER_S15_M5
`endif 

`ifdef AXI_AR_LAYER_S15_M6
  `undef AXI_AR_LAYER_S15_M6
`endif 

`ifdef AXI_AR_LAYER_S15_M7
  `undef AXI_AR_LAYER_S15_M7
`endif 

`ifdef AXI_AR_LAYER_S15_M8
  `undef AXI_AR_LAYER_S15_M8
`endif 

`ifdef AXI_AR_LAYER_S15_M9
  `undef AXI_AR_LAYER_S15_M9
`endif 

`ifdef AXI_AR_LAYER_S15_M10
  `undef AXI_AR_LAYER_S15_M10
`endif 

`ifdef AXI_AR_LAYER_S15_M11
  `undef AXI_AR_LAYER_S15_M11
`endif 

`ifdef AXI_AR_LAYER_S15_M12
  `undef AXI_AR_LAYER_S15_M12
`endif 

`ifdef AXI_AR_LAYER_S15_M13
  `undef AXI_AR_LAYER_S15_M13
`endif 

`ifdef AXI_AR_LAYER_S15_M14
  `undef AXI_AR_LAYER_S15_M14
`endif 

`ifdef AXI_AR_LAYER_S15_M15
  `undef AXI_AR_LAYER_S15_M15
`endif 

`ifdef AXI_AR_LAYER_S15_M16
  `undef AXI_AR_LAYER_S15_M16
`endif 

`ifdef AXI_AW_LAYER_S15_M1
  `undef AXI_AW_LAYER_S15_M1
`endif 

`ifdef AXI_AW_LAYER_S15_M2
  `undef AXI_AW_LAYER_S15_M2
`endif 

`ifdef AXI_AW_LAYER_S15_M3
  `undef AXI_AW_LAYER_S15_M3
`endif 

`ifdef AXI_AW_LAYER_S15_M4
  `undef AXI_AW_LAYER_S15_M4
`endif 

`ifdef AXI_AW_LAYER_S15_M5
  `undef AXI_AW_LAYER_S15_M5
`endif 

`ifdef AXI_AW_LAYER_S15_M6
  `undef AXI_AW_LAYER_S15_M6
`endif 

`ifdef AXI_AW_LAYER_S15_M7
  `undef AXI_AW_LAYER_S15_M7
`endif 

`ifdef AXI_AW_LAYER_S15_M8
  `undef AXI_AW_LAYER_S15_M8
`endif 

`ifdef AXI_AW_LAYER_S15_M9
  `undef AXI_AW_LAYER_S15_M9
`endif 

`ifdef AXI_AW_LAYER_S15_M10
  `undef AXI_AW_LAYER_S15_M10
`endif 

`ifdef AXI_AW_LAYER_S15_M11
  `undef AXI_AW_LAYER_S15_M11
`endif 

`ifdef AXI_AW_LAYER_S15_M12
  `undef AXI_AW_LAYER_S15_M12
`endif 

`ifdef AXI_AW_LAYER_S15_M13
  `undef AXI_AW_LAYER_S15_M13
`endif 

`ifdef AXI_AW_LAYER_S15_M14
  `undef AXI_AW_LAYER_S15_M14
`endif 

`ifdef AXI_AW_LAYER_S15_M15
  `undef AXI_AW_LAYER_S15_M15
`endif 

`ifdef AXI_AW_LAYER_S15_M16
  `undef AXI_AW_LAYER_S15_M16
`endif 

`ifdef AXI_W_LAYER_S15_M1
  `undef AXI_W_LAYER_S15_M1
`endif 

`ifdef AXI_W_LAYER_S15_M2
  `undef AXI_W_LAYER_S15_M2
`endif 

`ifdef AXI_W_LAYER_S15_M3
  `undef AXI_W_LAYER_S15_M3
`endif 

`ifdef AXI_W_LAYER_S15_M4
  `undef AXI_W_LAYER_S15_M4
`endif 

`ifdef AXI_W_LAYER_S15_M5
  `undef AXI_W_LAYER_S15_M5
`endif 

`ifdef AXI_W_LAYER_S15_M6
  `undef AXI_W_LAYER_S15_M6
`endif 

`ifdef AXI_W_LAYER_S15_M7
  `undef AXI_W_LAYER_S15_M7
`endif 

`ifdef AXI_W_LAYER_S15_M8
  `undef AXI_W_LAYER_S15_M8
`endif 

`ifdef AXI_W_LAYER_S15_M9
  `undef AXI_W_LAYER_S15_M9
`endif 

`ifdef AXI_W_LAYER_S15_M10
  `undef AXI_W_LAYER_S15_M10
`endif 

`ifdef AXI_W_LAYER_S15_M11
  `undef AXI_W_LAYER_S15_M11
`endif 

`ifdef AXI_W_LAYER_S15_M12
  `undef AXI_W_LAYER_S15_M12
`endif 

`ifdef AXI_W_LAYER_S15_M13
  `undef AXI_W_LAYER_S15_M13
`endif 

`ifdef AXI_W_LAYER_S15_M14
  `undef AXI_W_LAYER_S15_M14
`endif 

`ifdef AXI_W_LAYER_S15_M15
  `undef AXI_W_LAYER_S15_M15
`endif 

`ifdef AXI_W_LAYER_S15_M16
  `undef AXI_W_LAYER_S15_M16
`endif 

`ifdef AXI_AR_LAYER_S16_M1
  `undef AXI_AR_LAYER_S16_M1
`endif 

`ifdef AXI_AR_LAYER_S16_M2
  `undef AXI_AR_LAYER_S16_M2
`endif 

`ifdef AXI_AR_LAYER_S16_M3
  `undef AXI_AR_LAYER_S16_M3
`endif 

`ifdef AXI_AR_LAYER_S16_M4
  `undef AXI_AR_LAYER_S16_M4
`endif 

`ifdef AXI_AR_LAYER_S16_M5
  `undef AXI_AR_LAYER_S16_M5
`endif 

`ifdef AXI_AR_LAYER_S16_M6
  `undef AXI_AR_LAYER_S16_M6
`endif 

`ifdef AXI_AR_LAYER_S16_M7
  `undef AXI_AR_LAYER_S16_M7
`endif 

`ifdef AXI_AR_LAYER_S16_M8
  `undef AXI_AR_LAYER_S16_M8
`endif 

`ifdef AXI_AR_LAYER_S16_M9
  `undef AXI_AR_LAYER_S16_M9
`endif 

`ifdef AXI_AR_LAYER_S16_M10
  `undef AXI_AR_LAYER_S16_M10
`endif 

`ifdef AXI_AR_LAYER_S16_M11
  `undef AXI_AR_LAYER_S16_M11
`endif 

`ifdef AXI_AR_LAYER_S16_M12
  `undef AXI_AR_LAYER_S16_M12
`endif 

`ifdef AXI_AR_LAYER_S16_M13
  `undef AXI_AR_LAYER_S16_M13
`endif 

`ifdef AXI_AR_LAYER_S16_M14
  `undef AXI_AR_LAYER_S16_M14
`endif 

`ifdef AXI_AR_LAYER_S16_M15
  `undef AXI_AR_LAYER_S16_M15
`endif 

`ifdef AXI_AR_LAYER_S16_M16
  `undef AXI_AR_LAYER_S16_M16
`endif 

`ifdef AXI_AW_LAYER_S16_M1
  `undef AXI_AW_LAYER_S16_M1
`endif 

`ifdef AXI_AW_LAYER_S16_M2
  `undef AXI_AW_LAYER_S16_M2
`endif 

`ifdef AXI_AW_LAYER_S16_M3
  `undef AXI_AW_LAYER_S16_M3
`endif 

`ifdef AXI_AW_LAYER_S16_M4
  `undef AXI_AW_LAYER_S16_M4
`endif 

`ifdef AXI_AW_LAYER_S16_M5
  `undef AXI_AW_LAYER_S16_M5
`endif 

`ifdef AXI_AW_LAYER_S16_M6
  `undef AXI_AW_LAYER_S16_M6
`endif 

`ifdef AXI_AW_LAYER_S16_M7
  `undef AXI_AW_LAYER_S16_M7
`endif 

`ifdef AXI_AW_LAYER_S16_M8
  `undef AXI_AW_LAYER_S16_M8
`endif 

`ifdef AXI_AW_LAYER_S16_M9
  `undef AXI_AW_LAYER_S16_M9
`endif 

`ifdef AXI_AW_LAYER_S16_M10
  `undef AXI_AW_LAYER_S16_M10
`endif 

`ifdef AXI_AW_LAYER_S16_M11
  `undef AXI_AW_LAYER_S16_M11
`endif 

`ifdef AXI_AW_LAYER_S16_M12
  `undef AXI_AW_LAYER_S16_M12
`endif 

`ifdef AXI_AW_LAYER_S16_M13
  `undef AXI_AW_LAYER_S16_M13
`endif 

`ifdef AXI_AW_LAYER_S16_M14
  `undef AXI_AW_LAYER_S16_M14
`endif 

`ifdef AXI_AW_LAYER_S16_M15
  `undef AXI_AW_LAYER_S16_M15
`endif 

`ifdef AXI_AW_LAYER_S16_M16
  `undef AXI_AW_LAYER_S16_M16
`endif 

`ifdef AXI_W_LAYER_S16_M1
  `undef AXI_W_LAYER_S16_M1
`endif 

`ifdef AXI_W_LAYER_S16_M2
  `undef AXI_W_LAYER_S16_M2
`endif 

`ifdef AXI_W_LAYER_S16_M3
  `undef AXI_W_LAYER_S16_M3
`endif 

`ifdef AXI_W_LAYER_S16_M4
  `undef AXI_W_LAYER_S16_M4
`endif 

`ifdef AXI_W_LAYER_S16_M5
  `undef AXI_W_LAYER_S16_M5
`endif 

`ifdef AXI_W_LAYER_S16_M6
  `undef AXI_W_LAYER_S16_M6
`endif 

`ifdef AXI_W_LAYER_S16_M7
  `undef AXI_W_LAYER_S16_M7
`endif 

`ifdef AXI_W_LAYER_S16_M8
  `undef AXI_W_LAYER_S16_M8
`endif 

`ifdef AXI_W_LAYER_S16_M9
  `undef AXI_W_LAYER_S16_M9
`endif 

`ifdef AXI_W_LAYER_S16_M10
  `undef AXI_W_LAYER_S16_M10
`endif 

`ifdef AXI_W_LAYER_S16_M11
  `undef AXI_W_LAYER_S16_M11
`endif 

`ifdef AXI_W_LAYER_S16_M12
  `undef AXI_W_LAYER_S16_M12
`endif 

`ifdef AXI_W_LAYER_S16_M13
  `undef AXI_W_LAYER_S16_M13
`endif 

`ifdef AXI_W_LAYER_S16_M14
  `undef AXI_W_LAYER_S16_M14
`endif 

`ifdef AXI_W_LAYER_S16_M15
  `undef AXI_W_LAYER_S16_M15
`endif 

`ifdef AXI_W_LAYER_S16_M16
  `undef AXI_W_LAYER_S16_M16
`endif 

`ifdef AXI_ALL_R_LAYER_SHARED
  `undef AXI_ALL_R_LAYER_SHARED
`endif 

`ifdef AXI_R_LAYER_M1_S0
  `undef AXI_R_LAYER_M1_S0
`endif 

`ifdef AXI_R_LAYER_M1_S1
  `undef AXI_R_LAYER_M1_S1
`endif 

`ifdef AXI_R_LAYER_M1_S2
  `undef AXI_R_LAYER_M1_S2
`endif 

`ifdef AXI_R_LAYER_M1_S3
  `undef AXI_R_LAYER_M1_S3
`endif 

`ifdef AXI_R_LAYER_M1_S4
  `undef AXI_R_LAYER_M1_S4
`endif 

`ifdef AXI_R_LAYER_M1_S5
  `undef AXI_R_LAYER_M1_S5
`endif 

`ifdef AXI_R_LAYER_M1_S6
  `undef AXI_R_LAYER_M1_S6
`endif 

`ifdef AXI_R_LAYER_M1_S7
  `undef AXI_R_LAYER_M1_S7
`endif 

`ifdef AXI_R_LAYER_M1_S8
  `undef AXI_R_LAYER_M1_S8
`endif 

`ifdef AXI_R_LAYER_M1_S9
  `undef AXI_R_LAYER_M1_S9
`endif 

`ifdef AXI_R_LAYER_M1_S10
  `undef AXI_R_LAYER_M1_S10
`endif 

`ifdef AXI_R_LAYER_M1_S11
  `undef AXI_R_LAYER_M1_S11
`endif 

`ifdef AXI_R_LAYER_M1_S12
  `undef AXI_R_LAYER_M1_S12
`endif 

`ifdef AXI_R_LAYER_M1_S13
  `undef AXI_R_LAYER_M1_S13
`endif 

`ifdef AXI_R_LAYER_M1_S14
  `undef AXI_R_LAYER_M1_S14
`endif 

`ifdef AXI_R_LAYER_M1_S15
  `undef AXI_R_LAYER_M1_S15
`endif 

`ifdef AXI_R_LAYER_M1_S16
  `undef AXI_R_LAYER_M1_S16
`endif 

`ifdef AXI_ALL_B_LAYER_SHARED
  `undef AXI_ALL_B_LAYER_SHARED
`endif 

`ifdef AXI_B_LAYER_M1_S0
  `undef AXI_B_LAYER_M1_S0
`endif 

`ifdef AXI_B_LAYER_M1_S1
  `undef AXI_B_LAYER_M1_S1
`endif 

`ifdef AXI_B_LAYER_M1_S2
  `undef AXI_B_LAYER_M1_S2
`endif 

`ifdef AXI_B_LAYER_M1_S3
  `undef AXI_B_LAYER_M1_S3
`endif 

`ifdef AXI_B_LAYER_M1_S4
  `undef AXI_B_LAYER_M1_S4
`endif 

`ifdef AXI_B_LAYER_M1_S5
  `undef AXI_B_LAYER_M1_S5
`endif 

`ifdef AXI_B_LAYER_M1_S6
  `undef AXI_B_LAYER_M1_S6
`endif 

`ifdef AXI_B_LAYER_M1_S7
  `undef AXI_B_LAYER_M1_S7
`endif 

`ifdef AXI_B_LAYER_M1_S8
  `undef AXI_B_LAYER_M1_S8
`endif 

`ifdef AXI_B_LAYER_M1_S9
  `undef AXI_B_LAYER_M1_S9
`endif 

`ifdef AXI_B_LAYER_M1_S10
  `undef AXI_B_LAYER_M1_S10
`endif 

`ifdef AXI_B_LAYER_M1_S11
  `undef AXI_B_LAYER_M1_S11
`endif 

`ifdef AXI_B_LAYER_M1_S12
  `undef AXI_B_LAYER_M1_S12
`endif 

`ifdef AXI_B_LAYER_M1_S13
  `undef AXI_B_LAYER_M1_S13
`endif 

`ifdef AXI_B_LAYER_M1_S14
  `undef AXI_B_LAYER_M1_S14
`endif 

`ifdef AXI_B_LAYER_M1_S15
  `undef AXI_B_LAYER_M1_S15
`endif 

`ifdef AXI_B_LAYER_M1_S16
  `undef AXI_B_LAYER_M1_S16
`endif 

`ifdef AXI_R_LAYER_M2_S0
  `undef AXI_R_LAYER_M2_S0
`endif 

`ifdef AXI_R_LAYER_M2_S1
  `undef AXI_R_LAYER_M2_S1
`endif 

`ifdef AXI_R_LAYER_M2_S2
  `undef AXI_R_LAYER_M2_S2
`endif 

`ifdef AXI_R_LAYER_M2_S3
  `undef AXI_R_LAYER_M2_S3
`endif 

`ifdef AXI_R_LAYER_M2_S4
  `undef AXI_R_LAYER_M2_S4
`endif 

`ifdef AXI_R_LAYER_M2_S5
  `undef AXI_R_LAYER_M2_S5
`endif 

`ifdef AXI_R_LAYER_M2_S6
  `undef AXI_R_LAYER_M2_S6
`endif 

`ifdef AXI_R_LAYER_M2_S7
  `undef AXI_R_LAYER_M2_S7
`endif 

`ifdef AXI_R_LAYER_M2_S8
  `undef AXI_R_LAYER_M2_S8
`endif 

`ifdef AXI_R_LAYER_M2_S9
  `undef AXI_R_LAYER_M2_S9
`endif 

`ifdef AXI_R_LAYER_M2_S10
  `undef AXI_R_LAYER_M2_S10
`endif 

`ifdef AXI_R_LAYER_M2_S11
  `undef AXI_R_LAYER_M2_S11
`endif 

`ifdef AXI_R_LAYER_M2_S12
  `undef AXI_R_LAYER_M2_S12
`endif 

`ifdef AXI_R_LAYER_M2_S13
  `undef AXI_R_LAYER_M2_S13
`endif 

`ifdef AXI_R_LAYER_M2_S14
  `undef AXI_R_LAYER_M2_S14
`endif 

`ifdef AXI_R_LAYER_M2_S15
  `undef AXI_R_LAYER_M2_S15
`endif 

`ifdef AXI_R_LAYER_M2_S16
  `undef AXI_R_LAYER_M2_S16
`endif 

`ifdef AXI_B_LAYER_M2_S0
  `undef AXI_B_LAYER_M2_S0
`endif 

`ifdef AXI_B_LAYER_M2_S1
  `undef AXI_B_LAYER_M2_S1
`endif 

`ifdef AXI_B_LAYER_M2_S2
  `undef AXI_B_LAYER_M2_S2
`endif 

`ifdef AXI_B_LAYER_M2_S3
  `undef AXI_B_LAYER_M2_S3
`endif 

`ifdef AXI_B_LAYER_M2_S4
  `undef AXI_B_LAYER_M2_S4
`endif 

`ifdef AXI_B_LAYER_M2_S5
  `undef AXI_B_LAYER_M2_S5
`endif 

`ifdef AXI_B_LAYER_M2_S6
  `undef AXI_B_LAYER_M2_S6
`endif 

`ifdef AXI_B_LAYER_M2_S7
  `undef AXI_B_LAYER_M2_S7
`endif 

`ifdef AXI_B_LAYER_M2_S8
  `undef AXI_B_LAYER_M2_S8
`endif 

`ifdef AXI_B_LAYER_M2_S9
  `undef AXI_B_LAYER_M2_S9
`endif 

`ifdef AXI_B_LAYER_M2_S10
  `undef AXI_B_LAYER_M2_S10
`endif 

`ifdef AXI_B_LAYER_M2_S11
  `undef AXI_B_LAYER_M2_S11
`endif 

`ifdef AXI_B_LAYER_M2_S12
  `undef AXI_B_LAYER_M2_S12
`endif 

`ifdef AXI_B_LAYER_M2_S13
  `undef AXI_B_LAYER_M2_S13
`endif 

`ifdef AXI_B_LAYER_M2_S14
  `undef AXI_B_LAYER_M2_S14
`endif 

`ifdef AXI_B_LAYER_M2_S15
  `undef AXI_B_LAYER_M2_S15
`endif 

`ifdef AXI_B_LAYER_M2_S16
  `undef AXI_B_LAYER_M2_S16
`endif 

`ifdef AXI_R_LAYER_M3_S0
  `undef AXI_R_LAYER_M3_S0
`endif 

`ifdef AXI_R_LAYER_M3_S1
  `undef AXI_R_LAYER_M3_S1
`endif 

`ifdef AXI_R_LAYER_M3_S2
  `undef AXI_R_LAYER_M3_S2
`endif 

`ifdef AXI_R_LAYER_M3_S3
  `undef AXI_R_LAYER_M3_S3
`endif 

`ifdef AXI_R_LAYER_M3_S4
  `undef AXI_R_LAYER_M3_S4
`endif 

`ifdef AXI_R_LAYER_M3_S5
  `undef AXI_R_LAYER_M3_S5
`endif 

`ifdef AXI_R_LAYER_M3_S6
  `undef AXI_R_LAYER_M3_S6
`endif 

`ifdef AXI_R_LAYER_M3_S7
  `undef AXI_R_LAYER_M3_S7
`endif 

`ifdef AXI_R_LAYER_M3_S8
  `undef AXI_R_LAYER_M3_S8
`endif 

`ifdef AXI_R_LAYER_M3_S9
  `undef AXI_R_LAYER_M3_S9
`endif 

`ifdef AXI_R_LAYER_M3_S10
  `undef AXI_R_LAYER_M3_S10
`endif 

`ifdef AXI_R_LAYER_M3_S11
  `undef AXI_R_LAYER_M3_S11
`endif 

`ifdef AXI_R_LAYER_M3_S12
  `undef AXI_R_LAYER_M3_S12
`endif 

`ifdef AXI_R_LAYER_M3_S13
  `undef AXI_R_LAYER_M3_S13
`endif 

`ifdef AXI_R_LAYER_M3_S14
  `undef AXI_R_LAYER_M3_S14
`endif 

`ifdef AXI_R_LAYER_M3_S15
  `undef AXI_R_LAYER_M3_S15
`endif 

`ifdef AXI_R_LAYER_M3_S16
  `undef AXI_R_LAYER_M3_S16
`endif 

`ifdef AXI_B_LAYER_M3_S0
  `undef AXI_B_LAYER_M3_S0
`endif 

`ifdef AXI_B_LAYER_M3_S1
  `undef AXI_B_LAYER_M3_S1
`endif 

`ifdef AXI_B_LAYER_M3_S2
  `undef AXI_B_LAYER_M3_S2
`endif 

`ifdef AXI_B_LAYER_M3_S3
  `undef AXI_B_LAYER_M3_S3
`endif 

`ifdef AXI_B_LAYER_M3_S4
  `undef AXI_B_LAYER_M3_S4
`endif 

`ifdef AXI_B_LAYER_M3_S5
  `undef AXI_B_LAYER_M3_S5
`endif 

`ifdef AXI_B_LAYER_M3_S6
  `undef AXI_B_LAYER_M3_S6
`endif 

`ifdef AXI_B_LAYER_M3_S7
  `undef AXI_B_LAYER_M3_S7
`endif 

`ifdef AXI_B_LAYER_M3_S8
  `undef AXI_B_LAYER_M3_S8
`endif 

`ifdef AXI_B_LAYER_M3_S9
  `undef AXI_B_LAYER_M3_S9
`endif 

`ifdef AXI_B_LAYER_M3_S10
  `undef AXI_B_LAYER_M3_S10
`endif 

`ifdef AXI_B_LAYER_M3_S11
  `undef AXI_B_LAYER_M3_S11
`endif 

`ifdef AXI_B_LAYER_M3_S12
  `undef AXI_B_LAYER_M3_S12
`endif 

`ifdef AXI_B_LAYER_M3_S13
  `undef AXI_B_LAYER_M3_S13
`endif 

`ifdef AXI_B_LAYER_M3_S14
  `undef AXI_B_LAYER_M3_S14
`endif 

`ifdef AXI_B_LAYER_M3_S15
  `undef AXI_B_LAYER_M3_S15
`endif 

`ifdef AXI_B_LAYER_M3_S16
  `undef AXI_B_LAYER_M3_S16
`endif 

`ifdef AXI_R_LAYER_M4_S0
  `undef AXI_R_LAYER_M4_S0
`endif 

`ifdef AXI_R_LAYER_M4_S1
  `undef AXI_R_LAYER_M4_S1
`endif 

`ifdef AXI_R_LAYER_M4_S2
  `undef AXI_R_LAYER_M4_S2
`endif 

`ifdef AXI_R_LAYER_M4_S3
  `undef AXI_R_LAYER_M4_S3
`endif 

`ifdef AXI_R_LAYER_M4_S4
  `undef AXI_R_LAYER_M4_S4
`endif 

`ifdef AXI_R_LAYER_M4_S5
  `undef AXI_R_LAYER_M4_S5
`endif 

`ifdef AXI_R_LAYER_M4_S6
  `undef AXI_R_LAYER_M4_S6
`endif 

`ifdef AXI_R_LAYER_M4_S7
  `undef AXI_R_LAYER_M4_S7
`endif 

`ifdef AXI_R_LAYER_M4_S8
  `undef AXI_R_LAYER_M4_S8
`endif 

`ifdef AXI_R_LAYER_M4_S9
  `undef AXI_R_LAYER_M4_S9
`endif 

`ifdef AXI_R_LAYER_M4_S10
  `undef AXI_R_LAYER_M4_S10
`endif 

`ifdef AXI_R_LAYER_M4_S11
  `undef AXI_R_LAYER_M4_S11
`endif 

`ifdef AXI_R_LAYER_M4_S12
  `undef AXI_R_LAYER_M4_S12
`endif 

`ifdef AXI_R_LAYER_M4_S13
  `undef AXI_R_LAYER_M4_S13
`endif 

`ifdef AXI_R_LAYER_M4_S14
  `undef AXI_R_LAYER_M4_S14
`endif 

`ifdef AXI_R_LAYER_M4_S15
  `undef AXI_R_LAYER_M4_S15
`endif 

`ifdef AXI_R_LAYER_M4_S16
  `undef AXI_R_LAYER_M4_S16
`endif 

`ifdef AXI_B_LAYER_M4_S0
  `undef AXI_B_LAYER_M4_S0
`endif 

`ifdef AXI_B_LAYER_M4_S1
  `undef AXI_B_LAYER_M4_S1
`endif 

`ifdef AXI_B_LAYER_M4_S2
  `undef AXI_B_LAYER_M4_S2
`endif 

`ifdef AXI_B_LAYER_M4_S3
  `undef AXI_B_LAYER_M4_S3
`endif 

`ifdef AXI_B_LAYER_M4_S4
  `undef AXI_B_LAYER_M4_S4
`endif 

`ifdef AXI_B_LAYER_M4_S5
  `undef AXI_B_LAYER_M4_S5
`endif 

`ifdef AXI_B_LAYER_M4_S6
  `undef AXI_B_LAYER_M4_S6
`endif 

`ifdef AXI_B_LAYER_M4_S7
  `undef AXI_B_LAYER_M4_S7
`endif 

`ifdef AXI_B_LAYER_M4_S8
  `undef AXI_B_LAYER_M4_S8
`endif 

`ifdef AXI_B_LAYER_M4_S9
  `undef AXI_B_LAYER_M4_S9
`endif 

`ifdef AXI_B_LAYER_M4_S10
  `undef AXI_B_LAYER_M4_S10
`endif 

`ifdef AXI_B_LAYER_M4_S11
  `undef AXI_B_LAYER_M4_S11
`endif 

`ifdef AXI_B_LAYER_M4_S12
  `undef AXI_B_LAYER_M4_S12
`endif 

`ifdef AXI_B_LAYER_M4_S13
  `undef AXI_B_LAYER_M4_S13
`endif 

`ifdef AXI_B_LAYER_M4_S14
  `undef AXI_B_LAYER_M4_S14
`endif 

`ifdef AXI_B_LAYER_M4_S15
  `undef AXI_B_LAYER_M4_S15
`endif 

`ifdef AXI_B_LAYER_M4_S16
  `undef AXI_B_LAYER_M4_S16
`endif 

`ifdef AXI_R_LAYER_M5_S0
  `undef AXI_R_LAYER_M5_S0
`endif 

`ifdef AXI_R_LAYER_M5_S1
  `undef AXI_R_LAYER_M5_S1
`endif 

`ifdef AXI_R_LAYER_M5_S2
  `undef AXI_R_LAYER_M5_S2
`endif 

`ifdef AXI_R_LAYER_M5_S3
  `undef AXI_R_LAYER_M5_S3
`endif 

`ifdef AXI_R_LAYER_M5_S4
  `undef AXI_R_LAYER_M5_S4
`endif 

`ifdef AXI_R_LAYER_M5_S5
  `undef AXI_R_LAYER_M5_S5
`endif 

`ifdef AXI_R_LAYER_M5_S6
  `undef AXI_R_LAYER_M5_S6
`endif 

`ifdef AXI_R_LAYER_M5_S7
  `undef AXI_R_LAYER_M5_S7
`endif 

`ifdef AXI_R_LAYER_M5_S8
  `undef AXI_R_LAYER_M5_S8
`endif 

`ifdef AXI_R_LAYER_M5_S9
  `undef AXI_R_LAYER_M5_S9
`endif 

`ifdef AXI_R_LAYER_M5_S10
  `undef AXI_R_LAYER_M5_S10
`endif 

`ifdef AXI_R_LAYER_M5_S11
  `undef AXI_R_LAYER_M5_S11
`endif 

`ifdef AXI_R_LAYER_M5_S12
  `undef AXI_R_LAYER_M5_S12
`endif 

`ifdef AXI_R_LAYER_M5_S13
  `undef AXI_R_LAYER_M5_S13
`endif 

`ifdef AXI_R_LAYER_M5_S14
  `undef AXI_R_LAYER_M5_S14
`endif 

`ifdef AXI_R_LAYER_M5_S15
  `undef AXI_R_LAYER_M5_S15
`endif 

`ifdef AXI_R_LAYER_M5_S16
  `undef AXI_R_LAYER_M5_S16
`endif 

`ifdef AXI_B_LAYER_M5_S0
  `undef AXI_B_LAYER_M5_S0
`endif 

`ifdef AXI_B_LAYER_M5_S1
  `undef AXI_B_LAYER_M5_S1
`endif 

`ifdef AXI_B_LAYER_M5_S2
  `undef AXI_B_LAYER_M5_S2
`endif 

`ifdef AXI_B_LAYER_M5_S3
  `undef AXI_B_LAYER_M5_S3
`endif 

`ifdef AXI_B_LAYER_M5_S4
  `undef AXI_B_LAYER_M5_S4
`endif 

`ifdef AXI_B_LAYER_M5_S5
  `undef AXI_B_LAYER_M5_S5
`endif 

`ifdef AXI_B_LAYER_M5_S6
  `undef AXI_B_LAYER_M5_S6
`endif 

`ifdef AXI_B_LAYER_M5_S7
  `undef AXI_B_LAYER_M5_S7
`endif 

`ifdef AXI_B_LAYER_M5_S8
  `undef AXI_B_LAYER_M5_S8
`endif 

`ifdef AXI_B_LAYER_M5_S9
  `undef AXI_B_LAYER_M5_S9
`endif 

`ifdef AXI_B_LAYER_M5_S10
  `undef AXI_B_LAYER_M5_S10
`endif 

`ifdef AXI_B_LAYER_M5_S11
  `undef AXI_B_LAYER_M5_S11
`endif 

`ifdef AXI_B_LAYER_M5_S12
  `undef AXI_B_LAYER_M5_S12
`endif 

`ifdef AXI_B_LAYER_M5_S13
  `undef AXI_B_LAYER_M5_S13
`endif 

`ifdef AXI_B_LAYER_M5_S14
  `undef AXI_B_LAYER_M5_S14
`endif 

`ifdef AXI_B_LAYER_M5_S15
  `undef AXI_B_LAYER_M5_S15
`endif 

`ifdef AXI_B_LAYER_M5_S16
  `undef AXI_B_LAYER_M5_S16
`endif 

`ifdef AXI_R_LAYER_M6_S0
  `undef AXI_R_LAYER_M6_S0
`endif 

`ifdef AXI_R_LAYER_M6_S1
  `undef AXI_R_LAYER_M6_S1
`endif 

`ifdef AXI_R_LAYER_M6_S2
  `undef AXI_R_LAYER_M6_S2
`endif 

`ifdef AXI_R_LAYER_M6_S3
  `undef AXI_R_LAYER_M6_S3
`endif 

`ifdef AXI_R_LAYER_M6_S4
  `undef AXI_R_LAYER_M6_S4
`endif 

`ifdef AXI_R_LAYER_M6_S5
  `undef AXI_R_LAYER_M6_S5
`endif 

`ifdef AXI_R_LAYER_M6_S6
  `undef AXI_R_LAYER_M6_S6
`endif 

`ifdef AXI_R_LAYER_M6_S7
  `undef AXI_R_LAYER_M6_S7
`endif 

`ifdef AXI_R_LAYER_M6_S8
  `undef AXI_R_LAYER_M6_S8
`endif 

`ifdef AXI_R_LAYER_M6_S9
  `undef AXI_R_LAYER_M6_S9
`endif 

`ifdef AXI_R_LAYER_M6_S10
  `undef AXI_R_LAYER_M6_S10
`endif 

`ifdef AXI_R_LAYER_M6_S11
  `undef AXI_R_LAYER_M6_S11
`endif 

`ifdef AXI_R_LAYER_M6_S12
  `undef AXI_R_LAYER_M6_S12
`endif 

`ifdef AXI_R_LAYER_M6_S13
  `undef AXI_R_LAYER_M6_S13
`endif 

`ifdef AXI_R_LAYER_M6_S14
  `undef AXI_R_LAYER_M6_S14
`endif 

`ifdef AXI_R_LAYER_M6_S15
  `undef AXI_R_LAYER_M6_S15
`endif 

`ifdef AXI_R_LAYER_M6_S16
  `undef AXI_R_LAYER_M6_S16
`endif 

`ifdef AXI_B_LAYER_M6_S0
  `undef AXI_B_LAYER_M6_S0
`endif 

`ifdef AXI_B_LAYER_M6_S1
  `undef AXI_B_LAYER_M6_S1
`endif 

`ifdef AXI_B_LAYER_M6_S2
  `undef AXI_B_LAYER_M6_S2
`endif 

`ifdef AXI_B_LAYER_M6_S3
  `undef AXI_B_LAYER_M6_S3
`endif 

`ifdef AXI_B_LAYER_M6_S4
  `undef AXI_B_LAYER_M6_S4
`endif 

`ifdef AXI_B_LAYER_M6_S5
  `undef AXI_B_LAYER_M6_S5
`endif 

`ifdef AXI_B_LAYER_M6_S6
  `undef AXI_B_LAYER_M6_S6
`endif 

`ifdef AXI_B_LAYER_M6_S7
  `undef AXI_B_LAYER_M6_S7
`endif 

`ifdef AXI_B_LAYER_M6_S8
  `undef AXI_B_LAYER_M6_S8
`endif 

`ifdef AXI_B_LAYER_M6_S9
  `undef AXI_B_LAYER_M6_S9
`endif 

`ifdef AXI_B_LAYER_M6_S10
  `undef AXI_B_LAYER_M6_S10
`endif 

`ifdef AXI_B_LAYER_M6_S11
  `undef AXI_B_LAYER_M6_S11
`endif 

`ifdef AXI_B_LAYER_M6_S12
  `undef AXI_B_LAYER_M6_S12
`endif 

`ifdef AXI_B_LAYER_M6_S13
  `undef AXI_B_LAYER_M6_S13
`endif 

`ifdef AXI_B_LAYER_M6_S14
  `undef AXI_B_LAYER_M6_S14
`endif 

`ifdef AXI_B_LAYER_M6_S15
  `undef AXI_B_LAYER_M6_S15
`endif 

`ifdef AXI_B_LAYER_M6_S16
  `undef AXI_B_LAYER_M6_S16
`endif 

`ifdef AXI_R_LAYER_M7_S0
  `undef AXI_R_LAYER_M7_S0
`endif 

`ifdef AXI_R_LAYER_M7_S1
  `undef AXI_R_LAYER_M7_S1
`endif 

`ifdef AXI_R_LAYER_M7_S2
  `undef AXI_R_LAYER_M7_S2
`endif 

`ifdef AXI_R_LAYER_M7_S3
  `undef AXI_R_LAYER_M7_S3
`endif 

`ifdef AXI_R_LAYER_M7_S4
  `undef AXI_R_LAYER_M7_S4
`endif 

`ifdef AXI_R_LAYER_M7_S5
  `undef AXI_R_LAYER_M7_S5
`endif 

`ifdef AXI_R_LAYER_M7_S6
  `undef AXI_R_LAYER_M7_S6
`endif 

`ifdef AXI_R_LAYER_M7_S7
  `undef AXI_R_LAYER_M7_S7
`endif 

`ifdef AXI_R_LAYER_M7_S8
  `undef AXI_R_LAYER_M7_S8
`endif 

`ifdef AXI_R_LAYER_M7_S9
  `undef AXI_R_LAYER_M7_S9
`endif 

`ifdef AXI_R_LAYER_M7_S10
  `undef AXI_R_LAYER_M7_S10
`endif 

`ifdef AXI_R_LAYER_M7_S11
  `undef AXI_R_LAYER_M7_S11
`endif 

`ifdef AXI_R_LAYER_M7_S12
  `undef AXI_R_LAYER_M7_S12
`endif 

`ifdef AXI_R_LAYER_M7_S13
  `undef AXI_R_LAYER_M7_S13
`endif 

`ifdef AXI_R_LAYER_M7_S14
  `undef AXI_R_LAYER_M7_S14
`endif 

`ifdef AXI_R_LAYER_M7_S15
  `undef AXI_R_LAYER_M7_S15
`endif 

`ifdef AXI_R_LAYER_M7_S16
  `undef AXI_R_LAYER_M7_S16
`endif 

`ifdef AXI_B_LAYER_M7_S0
  `undef AXI_B_LAYER_M7_S0
`endif 

`ifdef AXI_B_LAYER_M7_S1
  `undef AXI_B_LAYER_M7_S1
`endif 

`ifdef AXI_B_LAYER_M7_S2
  `undef AXI_B_LAYER_M7_S2
`endif 

`ifdef AXI_B_LAYER_M7_S3
  `undef AXI_B_LAYER_M7_S3
`endif 

`ifdef AXI_B_LAYER_M7_S4
  `undef AXI_B_LAYER_M7_S4
`endif 

`ifdef AXI_B_LAYER_M7_S5
  `undef AXI_B_LAYER_M7_S5
`endif 

`ifdef AXI_B_LAYER_M7_S6
  `undef AXI_B_LAYER_M7_S6
`endif 

`ifdef AXI_B_LAYER_M7_S7
  `undef AXI_B_LAYER_M7_S7
`endif 

`ifdef AXI_B_LAYER_M7_S8
  `undef AXI_B_LAYER_M7_S8
`endif 

`ifdef AXI_B_LAYER_M7_S9
  `undef AXI_B_LAYER_M7_S9
`endif 

`ifdef AXI_B_LAYER_M7_S10
  `undef AXI_B_LAYER_M7_S10
`endif 

`ifdef AXI_B_LAYER_M7_S11
  `undef AXI_B_LAYER_M7_S11
`endif 

`ifdef AXI_B_LAYER_M7_S12
  `undef AXI_B_LAYER_M7_S12
`endif 

`ifdef AXI_B_LAYER_M7_S13
  `undef AXI_B_LAYER_M7_S13
`endif 

`ifdef AXI_B_LAYER_M7_S14
  `undef AXI_B_LAYER_M7_S14
`endif 

`ifdef AXI_B_LAYER_M7_S15
  `undef AXI_B_LAYER_M7_S15
`endif 

`ifdef AXI_B_LAYER_M7_S16
  `undef AXI_B_LAYER_M7_S16
`endif 

`ifdef AXI_R_LAYER_M8_S0
  `undef AXI_R_LAYER_M8_S0
`endif 

`ifdef AXI_R_LAYER_M8_S1
  `undef AXI_R_LAYER_M8_S1
`endif 

`ifdef AXI_R_LAYER_M8_S2
  `undef AXI_R_LAYER_M8_S2
`endif 

`ifdef AXI_R_LAYER_M8_S3
  `undef AXI_R_LAYER_M8_S3
`endif 

`ifdef AXI_R_LAYER_M8_S4
  `undef AXI_R_LAYER_M8_S4
`endif 

`ifdef AXI_R_LAYER_M8_S5
  `undef AXI_R_LAYER_M8_S5
`endif 

`ifdef AXI_R_LAYER_M8_S6
  `undef AXI_R_LAYER_M8_S6
`endif 

`ifdef AXI_R_LAYER_M8_S7
  `undef AXI_R_LAYER_M8_S7
`endif 

`ifdef AXI_R_LAYER_M8_S8
  `undef AXI_R_LAYER_M8_S8
`endif 

`ifdef AXI_R_LAYER_M8_S9
  `undef AXI_R_LAYER_M8_S9
`endif 

`ifdef AXI_R_LAYER_M8_S10
  `undef AXI_R_LAYER_M8_S10
`endif 

`ifdef AXI_R_LAYER_M8_S11
  `undef AXI_R_LAYER_M8_S11
`endif 

`ifdef AXI_R_LAYER_M8_S12
  `undef AXI_R_LAYER_M8_S12
`endif 

`ifdef AXI_R_LAYER_M8_S13
  `undef AXI_R_LAYER_M8_S13
`endif 

`ifdef AXI_R_LAYER_M8_S14
  `undef AXI_R_LAYER_M8_S14
`endif 

`ifdef AXI_R_LAYER_M8_S15
  `undef AXI_R_LAYER_M8_S15
`endif 

`ifdef AXI_R_LAYER_M8_S16
  `undef AXI_R_LAYER_M8_S16
`endif 

`ifdef AXI_B_LAYER_M8_S0
  `undef AXI_B_LAYER_M8_S0
`endif 

`ifdef AXI_B_LAYER_M8_S1
  `undef AXI_B_LAYER_M8_S1
`endif 

`ifdef AXI_B_LAYER_M8_S2
  `undef AXI_B_LAYER_M8_S2
`endif 

`ifdef AXI_B_LAYER_M8_S3
  `undef AXI_B_LAYER_M8_S3
`endif 

`ifdef AXI_B_LAYER_M8_S4
  `undef AXI_B_LAYER_M8_S4
`endif 

`ifdef AXI_B_LAYER_M8_S5
  `undef AXI_B_LAYER_M8_S5
`endif 

`ifdef AXI_B_LAYER_M8_S6
  `undef AXI_B_LAYER_M8_S6
`endif 

`ifdef AXI_B_LAYER_M8_S7
  `undef AXI_B_LAYER_M8_S7
`endif 

`ifdef AXI_B_LAYER_M8_S8
  `undef AXI_B_LAYER_M8_S8
`endif 

`ifdef AXI_B_LAYER_M8_S9
  `undef AXI_B_LAYER_M8_S9
`endif 

`ifdef AXI_B_LAYER_M8_S10
  `undef AXI_B_LAYER_M8_S10
`endif 

`ifdef AXI_B_LAYER_M8_S11
  `undef AXI_B_LAYER_M8_S11
`endif 

`ifdef AXI_B_LAYER_M8_S12
  `undef AXI_B_LAYER_M8_S12
`endif 

`ifdef AXI_B_LAYER_M8_S13
  `undef AXI_B_LAYER_M8_S13
`endif 

`ifdef AXI_B_LAYER_M8_S14
  `undef AXI_B_LAYER_M8_S14
`endif 

`ifdef AXI_B_LAYER_M8_S15
  `undef AXI_B_LAYER_M8_S15
`endif 

`ifdef AXI_B_LAYER_M8_S16
  `undef AXI_B_LAYER_M8_S16
`endif 

`ifdef AXI_R_LAYER_M9_S0
  `undef AXI_R_LAYER_M9_S0
`endif 

`ifdef AXI_R_LAYER_M9_S1
  `undef AXI_R_LAYER_M9_S1
`endif 

`ifdef AXI_R_LAYER_M9_S2
  `undef AXI_R_LAYER_M9_S2
`endif 

`ifdef AXI_R_LAYER_M9_S3
  `undef AXI_R_LAYER_M9_S3
`endif 

`ifdef AXI_R_LAYER_M9_S4
  `undef AXI_R_LAYER_M9_S4
`endif 

`ifdef AXI_R_LAYER_M9_S5
  `undef AXI_R_LAYER_M9_S5
`endif 

`ifdef AXI_R_LAYER_M9_S6
  `undef AXI_R_LAYER_M9_S6
`endif 

`ifdef AXI_R_LAYER_M9_S7
  `undef AXI_R_LAYER_M9_S7
`endif 

`ifdef AXI_R_LAYER_M9_S8
  `undef AXI_R_LAYER_M9_S8
`endif 

`ifdef AXI_R_LAYER_M9_S9
  `undef AXI_R_LAYER_M9_S9
`endif 

`ifdef AXI_R_LAYER_M9_S10
  `undef AXI_R_LAYER_M9_S10
`endif 

`ifdef AXI_R_LAYER_M9_S11
  `undef AXI_R_LAYER_M9_S11
`endif 

`ifdef AXI_R_LAYER_M9_S12
  `undef AXI_R_LAYER_M9_S12
`endif 

`ifdef AXI_R_LAYER_M9_S13
  `undef AXI_R_LAYER_M9_S13
`endif 

`ifdef AXI_R_LAYER_M9_S14
  `undef AXI_R_LAYER_M9_S14
`endif 

`ifdef AXI_R_LAYER_M9_S15
  `undef AXI_R_LAYER_M9_S15
`endif 

`ifdef AXI_R_LAYER_M9_S16
  `undef AXI_R_LAYER_M9_S16
`endif 

`ifdef AXI_B_LAYER_M9_S0
  `undef AXI_B_LAYER_M9_S0
`endif 

`ifdef AXI_B_LAYER_M9_S1
  `undef AXI_B_LAYER_M9_S1
`endif 

`ifdef AXI_B_LAYER_M9_S2
  `undef AXI_B_LAYER_M9_S2
`endif 

`ifdef AXI_B_LAYER_M9_S3
  `undef AXI_B_LAYER_M9_S3
`endif 

`ifdef AXI_B_LAYER_M9_S4
  `undef AXI_B_LAYER_M9_S4
`endif 

`ifdef AXI_B_LAYER_M9_S5
  `undef AXI_B_LAYER_M9_S5
`endif 

`ifdef AXI_B_LAYER_M9_S6
  `undef AXI_B_LAYER_M9_S6
`endif 

`ifdef AXI_B_LAYER_M9_S7
  `undef AXI_B_LAYER_M9_S7
`endif 

`ifdef AXI_B_LAYER_M9_S8
  `undef AXI_B_LAYER_M9_S8
`endif 

`ifdef AXI_B_LAYER_M9_S9
  `undef AXI_B_LAYER_M9_S9
`endif 

`ifdef AXI_B_LAYER_M9_S10
  `undef AXI_B_LAYER_M9_S10
`endif 

`ifdef AXI_B_LAYER_M9_S11
  `undef AXI_B_LAYER_M9_S11
`endif 

`ifdef AXI_B_LAYER_M9_S12
  `undef AXI_B_LAYER_M9_S12
`endif 

`ifdef AXI_B_LAYER_M9_S13
  `undef AXI_B_LAYER_M9_S13
`endif 

`ifdef AXI_B_LAYER_M9_S14
  `undef AXI_B_LAYER_M9_S14
`endif 

`ifdef AXI_B_LAYER_M9_S15
  `undef AXI_B_LAYER_M9_S15
`endif 

`ifdef AXI_B_LAYER_M9_S16
  `undef AXI_B_LAYER_M9_S16
`endif 

`ifdef AXI_R_LAYER_M10_S0
  `undef AXI_R_LAYER_M10_S0
`endif 

`ifdef AXI_R_LAYER_M10_S1
  `undef AXI_R_LAYER_M10_S1
`endif 

`ifdef AXI_R_LAYER_M10_S2
  `undef AXI_R_LAYER_M10_S2
`endif 

`ifdef AXI_R_LAYER_M10_S3
  `undef AXI_R_LAYER_M10_S3
`endif 

`ifdef AXI_R_LAYER_M10_S4
  `undef AXI_R_LAYER_M10_S4
`endif 

`ifdef AXI_R_LAYER_M10_S5
  `undef AXI_R_LAYER_M10_S5
`endif 

`ifdef AXI_R_LAYER_M10_S6
  `undef AXI_R_LAYER_M10_S6
`endif 

`ifdef AXI_R_LAYER_M10_S7
  `undef AXI_R_LAYER_M10_S7
`endif 

`ifdef AXI_R_LAYER_M10_S8
  `undef AXI_R_LAYER_M10_S8
`endif 

`ifdef AXI_R_LAYER_M10_S9
  `undef AXI_R_LAYER_M10_S9
`endif 

`ifdef AXI_R_LAYER_M10_S10
  `undef AXI_R_LAYER_M10_S10
`endif 

`ifdef AXI_R_LAYER_M10_S11
  `undef AXI_R_LAYER_M10_S11
`endif 

`ifdef AXI_R_LAYER_M10_S12
  `undef AXI_R_LAYER_M10_S12
`endif 

`ifdef AXI_R_LAYER_M10_S13
  `undef AXI_R_LAYER_M10_S13
`endif 

`ifdef AXI_R_LAYER_M10_S14
  `undef AXI_R_LAYER_M10_S14
`endif 

`ifdef AXI_R_LAYER_M10_S15
  `undef AXI_R_LAYER_M10_S15
`endif 

`ifdef AXI_R_LAYER_M10_S16
  `undef AXI_R_LAYER_M10_S16
`endif 

`ifdef AXI_B_LAYER_M10_S0
  `undef AXI_B_LAYER_M10_S0
`endif 

`ifdef AXI_B_LAYER_M10_S1
  `undef AXI_B_LAYER_M10_S1
`endif 

`ifdef AXI_B_LAYER_M10_S2
  `undef AXI_B_LAYER_M10_S2
`endif 

`ifdef AXI_B_LAYER_M10_S3
  `undef AXI_B_LAYER_M10_S3
`endif 

`ifdef AXI_B_LAYER_M10_S4
  `undef AXI_B_LAYER_M10_S4
`endif 

`ifdef AXI_B_LAYER_M10_S5
  `undef AXI_B_LAYER_M10_S5
`endif 

`ifdef AXI_B_LAYER_M10_S6
  `undef AXI_B_LAYER_M10_S6
`endif 

`ifdef AXI_B_LAYER_M10_S7
  `undef AXI_B_LAYER_M10_S7
`endif 

`ifdef AXI_B_LAYER_M10_S8
  `undef AXI_B_LAYER_M10_S8
`endif 

`ifdef AXI_B_LAYER_M10_S9
  `undef AXI_B_LAYER_M10_S9
`endif 

`ifdef AXI_B_LAYER_M10_S10
  `undef AXI_B_LAYER_M10_S10
`endif 

`ifdef AXI_B_LAYER_M10_S11
  `undef AXI_B_LAYER_M10_S11
`endif 

`ifdef AXI_B_LAYER_M10_S12
  `undef AXI_B_LAYER_M10_S12
`endif 

`ifdef AXI_B_LAYER_M10_S13
  `undef AXI_B_LAYER_M10_S13
`endif 

`ifdef AXI_B_LAYER_M10_S14
  `undef AXI_B_LAYER_M10_S14
`endif 

`ifdef AXI_B_LAYER_M10_S15
  `undef AXI_B_LAYER_M10_S15
`endif 

`ifdef AXI_B_LAYER_M10_S16
  `undef AXI_B_LAYER_M10_S16
`endif 

`ifdef AXI_R_LAYER_M11_S0
  `undef AXI_R_LAYER_M11_S0
`endif 

`ifdef AXI_R_LAYER_M11_S1
  `undef AXI_R_LAYER_M11_S1
`endif 

`ifdef AXI_R_LAYER_M11_S2
  `undef AXI_R_LAYER_M11_S2
`endif 

`ifdef AXI_R_LAYER_M11_S3
  `undef AXI_R_LAYER_M11_S3
`endif 

`ifdef AXI_R_LAYER_M11_S4
  `undef AXI_R_LAYER_M11_S4
`endif 

`ifdef AXI_R_LAYER_M11_S5
  `undef AXI_R_LAYER_M11_S5
`endif 

`ifdef AXI_R_LAYER_M11_S6
  `undef AXI_R_LAYER_M11_S6
`endif 

`ifdef AXI_R_LAYER_M11_S7
  `undef AXI_R_LAYER_M11_S7
`endif 

`ifdef AXI_R_LAYER_M11_S8
  `undef AXI_R_LAYER_M11_S8
`endif 

`ifdef AXI_R_LAYER_M11_S9
  `undef AXI_R_LAYER_M11_S9
`endif 

`ifdef AXI_R_LAYER_M11_S10
  `undef AXI_R_LAYER_M11_S10
`endif 

`ifdef AXI_R_LAYER_M11_S11
  `undef AXI_R_LAYER_M11_S11
`endif 

`ifdef AXI_R_LAYER_M11_S12
  `undef AXI_R_LAYER_M11_S12
`endif 

`ifdef AXI_R_LAYER_M11_S13
  `undef AXI_R_LAYER_M11_S13
`endif 

`ifdef AXI_R_LAYER_M11_S14
  `undef AXI_R_LAYER_M11_S14
`endif 

`ifdef AXI_R_LAYER_M11_S15
  `undef AXI_R_LAYER_M11_S15
`endif 

`ifdef AXI_R_LAYER_M11_S16
  `undef AXI_R_LAYER_M11_S16
`endif 

`ifdef AXI_B_LAYER_M11_S0
  `undef AXI_B_LAYER_M11_S0
`endif 

`ifdef AXI_B_LAYER_M11_S1
  `undef AXI_B_LAYER_M11_S1
`endif 

`ifdef AXI_B_LAYER_M11_S2
  `undef AXI_B_LAYER_M11_S2
`endif 

`ifdef AXI_B_LAYER_M11_S3
  `undef AXI_B_LAYER_M11_S3
`endif 

`ifdef AXI_B_LAYER_M11_S4
  `undef AXI_B_LAYER_M11_S4
`endif 

`ifdef AXI_B_LAYER_M11_S5
  `undef AXI_B_LAYER_M11_S5
`endif 

`ifdef AXI_B_LAYER_M11_S6
  `undef AXI_B_LAYER_M11_S6
`endif 

`ifdef AXI_B_LAYER_M11_S7
  `undef AXI_B_LAYER_M11_S7
`endif 

`ifdef AXI_B_LAYER_M11_S8
  `undef AXI_B_LAYER_M11_S8
`endif 

`ifdef AXI_B_LAYER_M11_S9
  `undef AXI_B_LAYER_M11_S9
`endif 

`ifdef AXI_B_LAYER_M11_S10
  `undef AXI_B_LAYER_M11_S10
`endif 

`ifdef AXI_B_LAYER_M11_S11
  `undef AXI_B_LAYER_M11_S11
`endif 

`ifdef AXI_B_LAYER_M11_S12
  `undef AXI_B_LAYER_M11_S12
`endif 

`ifdef AXI_B_LAYER_M11_S13
  `undef AXI_B_LAYER_M11_S13
`endif 

`ifdef AXI_B_LAYER_M11_S14
  `undef AXI_B_LAYER_M11_S14
`endif 

`ifdef AXI_B_LAYER_M11_S15
  `undef AXI_B_LAYER_M11_S15
`endif 

`ifdef AXI_B_LAYER_M11_S16
  `undef AXI_B_LAYER_M11_S16
`endif 

`ifdef AXI_R_LAYER_M12_S0
  `undef AXI_R_LAYER_M12_S0
`endif 

`ifdef AXI_R_LAYER_M12_S1
  `undef AXI_R_LAYER_M12_S1
`endif 

`ifdef AXI_R_LAYER_M12_S2
  `undef AXI_R_LAYER_M12_S2
`endif 

`ifdef AXI_R_LAYER_M12_S3
  `undef AXI_R_LAYER_M12_S3
`endif 

`ifdef AXI_R_LAYER_M12_S4
  `undef AXI_R_LAYER_M12_S4
`endif 

`ifdef AXI_R_LAYER_M12_S5
  `undef AXI_R_LAYER_M12_S5
`endif 

`ifdef AXI_R_LAYER_M12_S6
  `undef AXI_R_LAYER_M12_S6
`endif 

`ifdef AXI_R_LAYER_M12_S7
  `undef AXI_R_LAYER_M12_S7
`endif 

`ifdef AXI_R_LAYER_M12_S8
  `undef AXI_R_LAYER_M12_S8
`endif 

`ifdef AXI_R_LAYER_M12_S9
  `undef AXI_R_LAYER_M12_S9
`endif 

`ifdef AXI_R_LAYER_M12_S10
  `undef AXI_R_LAYER_M12_S10
`endif 

`ifdef AXI_R_LAYER_M12_S11
  `undef AXI_R_LAYER_M12_S11
`endif 

`ifdef AXI_R_LAYER_M12_S12
  `undef AXI_R_LAYER_M12_S12
`endif 

`ifdef AXI_R_LAYER_M12_S13
  `undef AXI_R_LAYER_M12_S13
`endif 

`ifdef AXI_R_LAYER_M12_S14
  `undef AXI_R_LAYER_M12_S14
`endif 

`ifdef AXI_R_LAYER_M12_S15
  `undef AXI_R_LAYER_M12_S15
`endif 

`ifdef AXI_R_LAYER_M12_S16
  `undef AXI_R_LAYER_M12_S16
`endif 

`ifdef AXI_B_LAYER_M12_S0
  `undef AXI_B_LAYER_M12_S0
`endif 

`ifdef AXI_B_LAYER_M12_S1
  `undef AXI_B_LAYER_M12_S1
`endif 

`ifdef AXI_B_LAYER_M12_S2
  `undef AXI_B_LAYER_M12_S2
`endif 

`ifdef AXI_B_LAYER_M12_S3
  `undef AXI_B_LAYER_M12_S3
`endif 

`ifdef AXI_B_LAYER_M12_S4
  `undef AXI_B_LAYER_M12_S4
`endif 

`ifdef AXI_B_LAYER_M12_S5
  `undef AXI_B_LAYER_M12_S5
`endif 

`ifdef AXI_B_LAYER_M12_S6
  `undef AXI_B_LAYER_M12_S6
`endif 

`ifdef AXI_B_LAYER_M12_S7
  `undef AXI_B_LAYER_M12_S7
`endif 

`ifdef AXI_B_LAYER_M12_S8
  `undef AXI_B_LAYER_M12_S8
`endif 

`ifdef AXI_B_LAYER_M12_S9
  `undef AXI_B_LAYER_M12_S9
`endif 

`ifdef AXI_B_LAYER_M12_S10
  `undef AXI_B_LAYER_M12_S10
`endif 

`ifdef AXI_B_LAYER_M12_S11
  `undef AXI_B_LAYER_M12_S11
`endif 

`ifdef AXI_B_LAYER_M12_S12
  `undef AXI_B_LAYER_M12_S12
`endif 

`ifdef AXI_B_LAYER_M12_S13
  `undef AXI_B_LAYER_M12_S13
`endif 

`ifdef AXI_B_LAYER_M12_S14
  `undef AXI_B_LAYER_M12_S14
`endif 

`ifdef AXI_B_LAYER_M12_S15
  `undef AXI_B_LAYER_M12_S15
`endif 

`ifdef AXI_B_LAYER_M12_S16
  `undef AXI_B_LAYER_M12_S16
`endif 

`ifdef AXI_R_LAYER_M13_S0
  `undef AXI_R_LAYER_M13_S0
`endif 

`ifdef AXI_R_LAYER_M13_S1
  `undef AXI_R_LAYER_M13_S1
`endif 

`ifdef AXI_R_LAYER_M13_S2
  `undef AXI_R_LAYER_M13_S2
`endif 

`ifdef AXI_R_LAYER_M13_S3
  `undef AXI_R_LAYER_M13_S3
`endif 

`ifdef AXI_R_LAYER_M13_S4
  `undef AXI_R_LAYER_M13_S4
`endif 

`ifdef AXI_R_LAYER_M13_S5
  `undef AXI_R_LAYER_M13_S5
`endif 

`ifdef AXI_R_LAYER_M13_S6
  `undef AXI_R_LAYER_M13_S6
`endif 

`ifdef AXI_R_LAYER_M13_S7
  `undef AXI_R_LAYER_M13_S7
`endif 

`ifdef AXI_R_LAYER_M13_S8
  `undef AXI_R_LAYER_M13_S8
`endif 

`ifdef AXI_R_LAYER_M13_S9
  `undef AXI_R_LAYER_M13_S9
`endif 

`ifdef AXI_R_LAYER_M13_S10
  `undef AXI_R_LAYER_M13_S10
`endif 

`ifdef AXI_R_LAYER_M13_S11
  `undef AXI_R_LAYER_M13_S11
`endif 

`ifdef AXI_R_LAYER_M13_S12
  `undef AXI_R_LAYER_M13_S12
`endif 

`ifdef AXI_R_LAYER_M13_S13
  `undef AXI_R_LAYER_M13_S13
`endif 

`ifdef AXI_R_LAYER_M13_S14
  `undef AXI_R_LAYER_M13_S14
`endif 

`ifdef AXI_R_LAYER_M13_S15
  `undef AXI_R_LAYER_M13_S15
`endif 

`ifdef AXI_R_LAYER_M13_S16
  `undef AXI_R_LAYER_M13_S16
`endif 

`ifdef AXI_B_LAYER_M13_S0
  `undef AXI_B_LAYER_M13_S0
`endif 

`ifdef AXI_B_LAYER_M13_S1
  `undef AXI_B_LAYER_M13_S1
`endif 

`ifdef AXI_B_LAYER_M13_S2
  `undef AXI_B_LAYER_M13_S2
`endif 

`ifdef AXI_B_LAYER_M13_S3
  `undef AXI_B_LAYER_M13_S3
`endif 

`ifdef AXI_B_LAYER_M13_S4
  `undef AXI_B_LAYER_M13_S4
`endif 

`ifdef AXI_B_LAYER_M13_S5
  `undef AXI_B_LAYER_M13_S5
`endif 

`ifdef AXI_B_LAYER_M13_S6
  `undef AXI_B_LAYER_M13_S6
`endif 

`ifdef AXI_B_LAYER_M13_S7
  `undef AXI_B_LAYER_M13_S7
`endif 

`ifdef AXI_B_LAYER_M13_S8
  `undef AXI_B_LAYER_M13_S8
`endif 

`ifdef AXI_B_LAYER_M13_S9
  `undef AXI_B_LAYER_M13_S9
`endif 

`ifdef AXI_B_LAYER_M13_S10
  `undef AXI_B_LAYER_M13_S10
`endif 

`ifdef AXI_B_LAYER_M13_S11
  `undef AXI_B_LAYER_M13_S11
`endif 

`ifdef AXI_B_LAYER_M13_S12
  `undef AXI_B_LAYER_M13_S12
`endif 

`ifdef AXI_B_LAYER_M13_S13
  `undef AXI_B_LAYER_M13_S13
`endif 

`ifdef AXI_B_LAYER_M13_S14
  `undef AXI_B_LAYER_M13_S14
`endif 

`ifdef AXI_B_LAYER_M13_S15
  `undef AXI_B_LAYER_M13_S15
`endif 

`ifdef AXI_B_LAYER_M13_S16
  `undef AXI_B_LAYER_M13_S16
`endif 

`ifdef AXI_R_LAYER_M14_S0
  `undef AXI_R_LAYER_M14_S0
`endif 

`ifdef AXI_R_LAYER_M14_S1
  `undef AXI_R_LAYER_M14_S1
`endif 

`ifdef AXI_R_LAYER_M14_S2
  `undef AXI_R_LAYER_M14_S2
`endif 

`ifdef AXI_R_LAYER_M14_S3
  `undef AXI_R_LAYER_M14_S3
`endif 

`ifdef AXI_R_LAYER_M14_S4
  `undef AXI_R_LAYER_M14_S4
`endif 

`ifdef AXI_R_LAYER_M14_S5
  `undef AXI_R_LAYER_M14_S5
`endif 

`ifdef AXI_R_LAYER_M14_S6
  `undef AXI_R_LAYER_M14_S6
`endif 

`ifdef AXI_R_LAYER_M14_S7
  `undef AXI_R_LAYER_M14_S7
`endif 

`ifdef AXI_R_LAYER_M14_S8
  `undef AXI_R_LAYER_M14_S8
`endif 

`ifdef AXI_R_LAYER_M14_S9
  `undef AXI_R_LAYER_M14_S9
`endif 

`ifdef AXI_R_LAYER_M14_S10
  `undef AXI_R_LAYER_M14_S10
`endif 

`ifdef AXI_R_LAYER_M14_S11
  `undef AXI_R_LAYER_M14_S11
`endif 

`ifdef AXI_R_LAYER_M14_S12
  `undef AXI_R_LAYER_M14_S12
`endif 

`ifdef AXI_R_LAYER_M14_S13
  `undef AXI_R_LAYER_M14_S13
`endif 

`ifdef AXI_R_LAYER_M14_S14
  `undef AXI_R_LAYER_M14_S14
`endif 

`ifdef AXI_R_LAYER_M14_S15
  `undef AXI_R_LAYER_M14_S15
`endif 

`ifdef AXI_R_LAYER_M14_S16
  `undef AXI_R_LAYER_M14_S16
`endif 

`ifdef AXI_B_LAYER_M14_S0
  `undef AXI_B_LAYER_M14_S0
`endif 

`ifdef AXI_B_LAYER_M14_S1
  `undef AXI_B_LAYER_M14_S1
`endif 

`ifdef AXI_B_LAYER_M14_S2
  `undef AXI_B_LAYER_M14_S2
`endif 

`ifdef AXI_B_LAYER_M14_S3
  `undef AXI_B_LAYER_M14_S3
`endif 

`ifdef AXI_B_LAYER_M14_S4
  `undef AXI_B_LAYER_M14_S4
`endif 

`ifdef AXI_B_LAYER_M14_S5
  `undef AXI_B_LAYER_M14_S5
`endif 

`ifdef AXI_B_LAYER_M14_S6
  `undef AXI_B_LAYER_M14_S6
`endif 

`ifdef AXI_B_LAYER_M14_S7
  `undef AXI_B_LAYER_M14_S7
`endif 

`ifdef AXI_B_LAYER_M14_S8
  `undef AXI_B_LAYER_M14_S8
`endif 

`ifdef AXI_B_LAYER_M14_S9
  `undef AXI_B_LAYER_M14_S9
`endif 

`ifdef AXI_B_LAYER_M14_S10
  `undef AXI_B_LAYER_M14_S10
`endif 

`ifdef AXI_B_LAYER_M14_S11
  `undef AXI_B_LAYER_M14_S11
`endif 

`ifdef AXI_B_LAYER_M14_S12
  `undef AXI_B_LAYER_M14_S12
`endif 

`ifdef AXI_B_LAYER_M14_S13
  `undef AXI_B_LAYER_M14_S13
`endif 

`ifdef AXI_B_LAYER_M14_S14
  `undef AXI_B_LAYER_M14_S14
`endif 

`ifdef AXI_B_LAYER_M14_S15
  `undef AXI_B_LAYER_M14_S15
`endif 

`ifdef AXI_B_LAYER_M14_S16
  `undef AXI_B_LAYER_M14_S16
`endif 

`ifdef AXI_R_LAYER_M15_S0
  `undef AXI_R_LAYER_M15_S0
`endif 

`ifdef AXI_R_LAYER_M15_S1
  `undef AXI_R_LAYER_M15_S1
`endif 

`ifdef AXI_R_LAYER_M15_S2
  `undef AXI_R_LAYER_M15_S2
`endif 

`ifdef AXI_R_LAYER_M15_S3
  `undef AXI_R_LAYER_M15_S3
`endif 

`ifdef AXI_R_LAYER_M15_S4
  `undef AXI_R_LAYER_M15_S4
`endif 

`ifdef AXI_R_LAYER_M15_S5
  `undef AXI_R_LAYER_M15_S5
`endif 

`ifdef AXI_R_LAYER_M15_S6
  `undef AXI_R_LAYER_M15_S6
`endif 

`ifdef AXI_R_LAYER_M15_S7
  `undef AXI_R_LAYER_M15_S7
`endif 

`ifdef AXI_R_LAYER_M15_S8
  `undef AXI_R_LAYER_M15_S8
`endif 

`ifdef AXI_R_LAYER_M15_S9
  `undef AXI_R_LAYER_M15_S9
`endif 

`ifdef AXI_R_LAYER_M15_S10
  `undef AXI_R_LAYER_M15_S10
`endif 

`ifdef AXI_R_LAYER_M15_S11
  `undef AXI_R_LAYER_M15_S11
`endif 

`ifdef AXI_R_LAYER_M15_S12
  `undef AXI_R_LAYER_M15_S12
`endif 

`ifdef AXI_R_LAYER_M15_S13
  `undef AXI_R_LAYER_M15_S13
`endif 

`ifdef AXI_R_LAYER_M15_S14
  `undef AXI_R_LAYER_M15_S14
`endif 

`ifdef AXI_R_LAYER_M15_S15
  `undef AXI_R_LAYER_M15_S15
`endif 

`ifdef AXI_R_LAYER_M15_S16
  `undef AXI_R_LAYER_M15_S16
`endif 

`ifdef AXI_B_LAYER_M15_S0
  `undef AXI_B_LAYER_M15_S0
`endif 

`ifdef AXI_B_LAYER_M15_S1
  `undef AXI_B_LAYER_M15_S1
`endif 

`ifdef AXI_B_LAYER_M15_S2
  `undef AXI_B_LAYER_M15_S2
`endif 

`ifdef AXI_B_LAYER_M15_S3
  `undef AXI_B_LAYER_M15_S3
`endif 

`ifdef AXI_B_LAYER_M15_S4
  `undef AXI_B_LAYER_M15_S4
`endif 

`ifdef AXI_B_LAYER_M15_S5
  `undef AXI_B_LAYER_M15_S5
`endif 

`ifdef AXI_B_LAYER_M15_S6
  `undef AXI_B_LAYER_M15_S6
`endif 

`ifdef AXI_B_LAYER_M15_S7
  `undef AXI_B_LAYER_M15_S7
`endif 

`ifdef AXI_B_LAYER_M15_S8
  `undef AXI_B_LAYER_M15_S8
`endif 

`ifdef AXI_B_LAYER_M15_S9
  `undef AXI_B_LAYER_M15_S9
`endif 

`ifdef AXI_B_LAYER_M15_S10
  `undef AXI_B_LAYER_M15_S10
`endif 

`ifdef AXI_B_LAYER_M15_S11
  `undef AXI_B_LAYER_M15_S11
`endif 

`ifdef AXI_B_LAYER_M15_S12
  `undef AXI_B_LAYER_M15_S12
`endif 

`ifdef AXI_B_LAYER_M15_S13
  `undef AXI_B_LAYER_M15_S13
`endif 

`ifdef AXI_B_LAYER_M15_S14
  `undef AXI_B_LAYER_M15_S14
`endif 

`ifdef AXI_B_LAYER_M15_S15
  `undef AXI_B_LAYER_M15_S15
`endif 

`ifdef AXI_B_LAYER_M15_S16
  `undef AXI_B_LAYER_M15_S16
`endif 

`ifdef AXI_R_LAYER_M16_S0
  `undef AXI_R_LAYER_M16_S0
`endif 

`ifdef AXI_R_LAYER_M16_S1
  `undef AXI_R_LAYER_M16_S1
`endif 

`ifdef AXI_R_LAYER_M16_S2
  `undef AXI_R_LAYER_M16_S2
`endif 

`ifdef AXI_R_LAYER_M16_S3
  `undef AXI_R_LAYER_M16_S3
`endif 

`ifdef AXI_R_LAYER_M16_S4
  `undef AXI_R_LAYER_M16_S4
`endif 

`ifdef AXI_R_LAYER_M16_S5
  `undef AXI_R_LAYER_M16_S5
`endif 

`ifdef AXI_R_LAYER_M16_S6
  `undef AXI_R_LAYER_M16_S6
`endif 

`ifdef AXI_R_LAYER_M16_S7
  `undef AXI_R_LAYER_M16_S7
`endif 

`ifdef AXI_R_LAYER_M16_S8
  `undef AXI_R_LAYER_M16_S8
`endif 

`ifdef AXI_R_LAYER_M16_S9
  `undef AXI_R_LAYER_M16_S9
`endif 

`ifdef AXI_R_LAYER_M16_S10
  `undef AXI_R_LAYER_M16_S10
`endif 

`ifdef AXI_R_LAYER_M16_S11
  `undef AXI_R_LAYER_M16_S11
`endif 

`ifdef AXI_R_LAYER_M16_S12
  `undef AXI_R_LAYER_M16_S12
`endif 

`ifdef AXI_R_LAYER_M16_S13
  `undef AXI_R_LAYER_M16_S13
`endif 

`ifdef AXI_R_LAYER_M16_S14
  `undef AXI_R_LAYER_M16_S14
`endif 

`ifdef AXI_R_LAYER_M16_S15
  `undef AXI_R_LAYER_M16_S15
`endif 

`ifdef AXI_R_LAYER_M16_S16
  `undef AXI_R_LAYER_M16_S16
`endif 

`ifdef AXI_B_LAYER_M16_S0
  `undef AXI_B_LAYER_M16_S0
`endif 

`ifdef AXI_B_LAYER_M16_S1
  `undef AXI_B_LAYER_M16_S1
`endif 

`ifdef AXI_B_LAYER_M16_S2
  `undef AXI_B_LAYER_M16_S2
`endif 

`ifdef AXI_B_LAYER_M16_S3
  `undef AXI_B_LAYER_M16_S3
`endif 

`ifdef AXI_B_LAYER_M16_S4
  `undef AXI_B_LAYER_M16_S4
`endif 

`ifdef AXI_B_LAYER_M16_S5
  `undef AXI_B_LAYER_M16_S5
`endif 

`ifdef AXI_B_LAYER_M16_S6
  `undef AXI_B_LAYER_M16_S6
`endif 

`ifdef AXI_B_LAYER_M16_S7
  `undef AXI_B_LAYER_M16_S7
`endif 

`ifdef AXI_B_LAYER_M16_S8
  `undef AXI_B_LAYER_M16_S8
`endif 

`ifdef AXI_B_LAYER_M16_S9
  `undef AXI_B_LAYER_M16_S9
`endif 

`ifdef AXI_B_LAYER_M16_S10
  `undef AXI_B_LAYER_M16_S10
`endif 

`ifdef AXI_B_LAYER_M16_S11
  `undef AXI_B_LAYER_M16_S11
`endif 

`ifdef AXI_B_LAYER_M16_S12
  `undef AXI_B_LAYER_M16_S12
`endif 

`ifdef AXI_B_LAYER_M16_S13
  `undef AXI_B_LAYER_M16_S13
`endif 

`ifdef AXI_B_LAYER_M16_S14
  `undef AXI_B_LAYER_M16_S14
`endif 

`ifdef AXI_B_LAYER_M16_S15
  `undef AXI_B_LAYER_M16_S15
`endif 

`ifdef AXI_B_LAYER_M16_S16
  `undef AXI_B_LAYER_M16_S16
`endif 

`ifdef AXI_AR_HAS_SHARED_LAYER
  `undef AXI_AR_HAS_SHARED_LAYER
`endif 

`ifdef AXI_AR_SHARED_LAYER
  `undef AXI_AR_SHARED_LAYER
`endif 

`ifdef AXI_AW_HAS_SHARED_LAYER
  `undef AXI_AW_HAS_SHARED_LAYER
`endif 

`ifdef AXI_AW_SHARED_LAYER
  `undef AXI_AW_SHARED_LAYER
`endif 

`ifdef AXI_W_HAS_SHARED_LAYER
  `undef AXI_W_HAS_SHARED_LAYER
`endif 

`ifdef AXI_W_SHARED_LAYER
  `undef AXI_W_SHARED_LAYER
`endif 

`ifdef AXI_R_HAS_SHARED_LAYER
  `undef AXI_R_HAS_SHARED_LAYER
`endif 

`ifdef AXI_R_SHARED_LAYER
  `undef AXI_R_SHARED_LAYER
`endif 

`ifdef AXI_B_HAS_SHARED_LAYER
  `undef AXI_B_HAS_SHARED_LAYER
`endif 

`ifdef AXI_B_SHARED_LAYER
  `undef AXI_B_SHARED_LAYER
`endif 

`ifdef AXI_AR_SHARED_LAYER_NM
  `undef AXI_AR_SHARED_LAYER_NM
`endif 

`ifdef AXI_LOG2_AR_SHARED_LAYER_NM
  `undef AXI_LOG2_AR_SHARED_LAYER_NM
`endif 

`ifdef AXI_LOG2_AR_SHARED_LAYER_NMP1
  `undef AXI_LOG2_AR_SHARED_LAYER_NMP1
`endif 

`ifdef AXI_AR_SHARED_LAYER_NS
  `undef AXI_AR_SHARED_LAYER_NS
`endif 

`ifdef AXI_AR_SHARED_LAYER_NS_R0
  `undef AXI_AR_SHARED_LAYER_NS_R0
`endif 

`ifdef AXI_LOG2_AR_SHARED_LAYER_NS
  `undef AXI_LOG2_AR_SHARED_LAYER_NS
`endif 

`ifdef AXI_LOG2_AR_SHARED_LAYER_NSP1
  `undef AXI_LOG2_AR_SHARED_LAYER_NSP1
`endif 

`ifdef AXI_AW_SHARED_LAYER_NM
  `undef AXI_AW_SHARED_LAYER_NM
`endif 

`ifdef AXI_LOG2_AW_SHARED_LAYER_NM
  `undef AXI_LOG2_AW_SHARED_LAYER_NM
`endif 

`ifdef AXI_LOG2_AW_SHARED_LAYER_NMP1
  `undef AXI_LOG2_AW_SHARED_LAYER_NMP1
`endif 

`ifdef AXI_AW_SHARED_LAYER_NS
  `undef AXI_AW_SHARED_LAYER_NS
`endif 

`ifdef AXI_AW_SHARED_LAYER_NS_R0
  `undef AXI_AW_SHARED_LAYER_NS_R0
`endif 

`ifdef AXI_LOG2_AW_SHARED_LAYER_NS
  `undef AXI_LOG2_AW_SHARED_LAYER_NS
`endif 

`ifdef AXI_LOG2_AW_SHARED_LAYER_NSP1
  `undef AXI_LOG2_AW_SHARED_LAYER_NSP1
`endif 

`ifdef AXI_W_SHARED_LAYER_NM
  `undef AXI_W_SHARED_LAYER_NM
`endif 

`ifdef AXI_LOG2_W_SHARED_LAYER_NM
  `undef AXI_LOG2_W_SHARED_LAYER_NM
`endif 

`ifdef AXI_LOG2_W_SHARED_LAYER_NMP1
  `undef AXI_LOG2_W_SHARED_LAYER_NMP1
`endif 

`ifdef AXI_W_SHARED_LAYER_NS
  `undef AXI_W_SHARED_LAYER_NS
`endif 

`ifdef AXI_W_SHARED_LAYER_NS_R0
  `undef AXI_W_SHARED_LAYER_NS_R0
`endif 

`ifdef AXI_LOG2_W_SHARED_LAYER_NS
  `undef AXI_LOG2_W_SHARED_LAYER_NS
`endif 

`ifdef AXI_LOG2_W_SHARED_LAYER_NSP1
  `undef AXI_LOG2_W_SHARED_LAYER_NSP1
`endif 

`ifdef AXI_R_SHARED_LAYER_NM
  `undef AXI_R_SHARED_LAYER_NM
`endif 

`ifdef AXI_R_SHARED_LAYER_NM_R0
  `undef AXI_R_SHARED_LAYER_NM_R0
`endif 

`ifdef AXI_LOG2_R_SHARED_LAYER_NM
  `undef AXI_LOG2_R_SHARED_LAYER_NM
`endif 

`ifdef AXI_LOG2_R_SHARED_LAYER_NMP1
  `undef AXI_LOG2_R_SHARED_LAYER_NMP1
`endif 

`ifdef AXI_R_SHARED_LAYER_NS
  `undef AXI_R_SHARED_LAYER_NS
`endif 

`ifdef AXI_LOG2_R_SHARED_LAYER_NS
  `undef AXI_LOG2_R_SHARED_LAYER_NS
`endif 

`ifdef AXI_LOG2_R_SHARED_LAYER_NSP1
  `undef AXI_LOG2_R_SHARED_LAYER_NSP1
`endif 

`ifdef AXI_B_SHARED_LAYER_NM
  `undef AXI_B_SHARED_LAYER_NM
`endif 

`ifdef AXI_B_SHARED_LAYER_NM_R0
  `undef AXI_B_SHARED_LAYER_NM_R0
`endif 

`ifdef AXI_LOG2_B_SHARED_LAYER_NM
  `undef AXI_LOG2_B_SHARED_LAYER_NM
`endif 

`ifdef AXI_LOG2_B_SHARED_LAYER_NMP1
  `undef AXI_LOG2_B_SHARED_LAYER_NMP1
`endif 

`ifdef AXI_B_SHARED_LAYER_NS
  `undef AXI_B_SHARED_LAYER_NS
`endif 

`ifdef AXI_LOG2_B_SHARED_LAYER_NS
  `undef AXI_LOG2_B_SHARED_LAYER_NS
`endif 

`ifdef AXI_LOG2_B_SHARED_LAYER_NSP1
  `undef AXI_LOG2_B_SHARED_LAYER_NSP1
`endif 

`ifdef AXI_AR_S0_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AR_S0_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AR_S0_HAS_SHRD_DDCTD_LNK
  `undef AXI_AR_S0_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AR_S0_NMV
  `undef AXI_AR_S0_NMV
`endif 

`ifdef AXI_AR_S0_NMV_LOG2
  `undef AXI_AR_S0_NMV_LOG2
`endif 

`ifdef AXI_AR_S0_NMV_P1_LOG2
  `undef AXI_AR_S0_NMV_P1_LOG2
`endif 

`ifdef AXI_AW_S0_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AW_S0_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AW_S0_HAS_SHRD_DDCTD_LNK
  `undef AXI_AW_S0_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AW_S0_NMV
  `undef AXI_AW_S0_NMV
`endif 

`ifdef AXI_AW_S0_NMV_LOG2
  `undef AXI_AW_S0_NMV_LOG2
`endif 

`ifdef AXI_AW_S0_NMV_P1_LOG2
  `undef AXI_AW_S0_NMV_P1_LOG2
`endif 

`ifdef AXI_W_S0_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_W_S0_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_W_S0_HAS_SHRD_DDCTD_LNK
  `undef AXI_W_S0_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_W_S0_NMV
  `undef AXI_W_S0_NMV
`endif 

`ifdef AXI_W_S0_NMV_LOG2
  `undef AXI_W_S0_NMV_LOG2
`endif 

`ifdef AXI_W_S0_NMV_P1_LOG2
  `undef AXI_W_S0_NMV_P1_LOG2
`endif 

`ifdef AXI_AR_S1_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AR_S1_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AR_S1_HAS_SHRD_DDCTD_LNK
  `undef AXI_AR_S1_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AR_S1_NMV
  `undef AXI_AR_S1_NMV
`endif 

`ifdef AXI_AR_S1_NMV_LOG2
  `undef AXI_AR_S1_NMV_LOG2
`endif 

`ifdef AXI_AR_S1_NMV_P1_LOG2
  `undef AXI_AR_S1_NMV_P1_LOG2
`endif 

`ifdef AXI_AW_S1_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AW_S1_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AW_S1_HAS_SHRD_DDCTD_LNK
  `undef AXI_AW_S1_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AW_S1_NMV
  `undef AXI_AW_S1_NMV
`endif 

`ifdef AXI_AW_S1_NMV_LOG2
  `undef AXI_AW_S1_NMV_LOG2
`endif 

`ifdef AXI_AW_S1_NMV_P1_LOG2
  `undef AXI_AW_S1_NMV_P1_LOG2
`endif 

`ifdef AXI_W_S1_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_W_S1_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_W_S1_HAS_SHRD_DDCTD_LNK
  `undef AXI_W_S1_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_W_S1_NMV
  `undef AXI_W_S1_NMV
`endif 

`ifdef AXI_W_S1_NMV_LOG2
  `undef AXI_W_S1_NMV_LOG2
`endif 

`ifdef AXI_W_S1_NMV_P1_LOG2
  `undef AXI_W_S1_NMV_P1_LOG2
`endif 

`ifdef AXI_AR_S2_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AR_S2_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AR_S2_HAS_SHRD_DDCTD_LNK
  `undef AXI_AR_S2_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AR_S2_NMV
  `undef AXI_AR_S2_NMV
`endif 

`ifdef AXI_AR_S2_NMV_LOG2
  `undef AXI_AR_S2_NMV_LOG2
`endif 

`ifdef AXI_AR_S2_NMV_P1_LOG2
  `undef AXI_AR_S2_NMV_P1_LOG2
`endif 

`ifdef AXI_AW_S2_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AW_S2_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AW_S2_HAS_SHRD_DDCTD_LNK
  `undef AXI_AW_S2_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AW_S2_NMV
  `undef AXI_AW_S2_NMV
`endif 

`ifdef AXI_AW_S2_NMV_LOG2
  `undef AXI_AW_S2_NMV_LOG2
`endif 

`ifdef AXI_AW_S2_NMV_P1_LOG2
  `undef AXI_AW_S2_NMV_P1_LOG2
`endif 

`ifdef AXI_W_S2_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_W_S2_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_W_S2_HAS_SHRD_DDCTD_LNK
  `undef AXI_W_S2_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_W_S2_NMV
  `undef AXI_W_S2_NMV
`endif 

`ifdef AXI_W_S2_NMV_LOG2
  `undef AXI_W_S2_NMV_LOG2
`endif 

`ifdef AXI_W_S2_NMV_P1_LOG2
  `undef AXI_W_S2_NMV_P1_LOG2
`endif 

`ifdef AXI_AR_S3_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AR_S3_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AR_S3_HAS_SHRD_DDCTD_LNK
  `undef AXI_AR_S3_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AR_S3_NMV
  `undef AXI_AR_S3_NMV
`endif 

`ifdef AXI_AR_S3_NMV_LOG2
  `undef AXI_AR_S3_NMV_LOG2
`endif 

`ifdef AXI_AR_S3_NMV_P1_LOG2
  `undef AXI_AR_S3_NMV_P1_LOG2
`endif 

`ifdef AXI_AW_S3_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AW_S3_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AW_S3_HAS_SHRD_DDCTD_LNK
  `undef AXI_AW_S3_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AW_S3_NMV
  `undef AXI_AW_S3_NMV
`endif 

`ifdef AXI_AW_S3_NMV_LOG2
  `undef AXI_AW_S3_NMV_LOG2
`endif 

`ifdef AXI_AW_S3_NMV_P1_LOG2
  `undef AXI_AW_S3_NMV_P1_LOG2
`endif 

`ifdef AXI_W_S3_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_W_S3_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_W_S3_HAS_SHRD_DDCTD_LNK
  `undef AXI_W_S3_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_W_S3_NMV
  `undef AXI_W_S3_NMV
`endif 

`ifdef AXI_W_S3_NMV_LOG2
  `undef AXI_W_S3_NMV_LOG2
`endif 

`ifdef AXI_W_S3_NMV_P1_LOG2
  `undef AXI_W_S3_NMV_P1_LOG2
`endif 

`ifdef AXI_AR_S4_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AR_S4_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AR_S4_HAS_SHRD_DDCTD_LNK
  `undef AXI_AR_S4_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AR_S4_NMV
  `undef AXI_AR_S4_NMV
`endif 

`ifdef AXI_AR_S4_NMV_LOG2
  `undef AXI_AR_S4_NMV_LOG2
`endif 

`ifdef AXI_AR_S4_NMV_P1_LOG2
  `undef AXI_AR_S4_NMV_P1_LOG2
`endif 

`ifdef AXI_AW_S4_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AW_S4_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AW_S4_HAS_SHRD_DDCTD_LNK
  `undef AXI_AW_S4_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AW_S4_NMV
  `undef AXI_AW_S4_NMV
`endif 

`ifdef AXI_AW_S4_NMV_LOG2
  `undef AXI_AW_S4_NMV_LOG2
`endif 

`ifdef AXI_AW_S4_NMV_P1_LOG2
  `undef AXI_AW_S4_NMV_P1_LOG2
`endif 

`ifdef AXI_W_S4_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_W_S4_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_W_S4_HAS_SHRD_DDCTD_LNK
  `undef AXI_W_S4_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_W_S4_NMV
  `undef AXI_W_S4_NMV
`endif 

`ifdef AXI_W_S4_NMV_LOG2
  `undef AXI_W_S4_NMV_LOG2
`endif 

`ifdef AXI_W_S4_NMV_P1_LOG2
  `undef AXI_W_S4_NMV_P1_LOG2
`endif 

`ifdef AXI_AR_S5_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AR_S5_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AR_S5_HAS_SHRD_DDCTD_LNK
  `undef AXI_AR_S5_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AR_S5_NMV
  `undef AXI_AR_S5_NMV
`endif 

`ifdef AXI_AR_S5_NMV_LOG2
  `undef AXI_AR_S5_NMV_LOG2
`endif 

`ifdef AXI_AR_S5_NMV_P1_LOG2
  `undef AXI_AR_S5_NMV_P1_LOG2
`endif 

`ifdef AXI_AW_S5_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AW_S5_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AW_S5_HAS_SHRD_DDCTD_LNK
  `undef AXI_AW_S5_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AW_S5_NMV
  `undef AXI_AW_S5_NMV
`endif 

`ifdef AXI_AW_S5_NMV_LOG2
  `undef AXI_AW_S5_NMV_LOG2
`endif 

`ifdef AXI_AW_S5_NMV_P1_LOG2
  `undef AXI_AW_S5_NMV_P1_LOG2
`endif 

`ifdef AXI_W_S5_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_W_S5_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_W_S5_HAS_SHRD_DDCTD_LNK
  `undef AXI_W_S5_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_W_S5_NMV
  `undef AXI_W_S5_NMV
`endif 

`ifdef AXI_W_S5_NMV_LOG2
  `undef AXI_W_S5_NMV_LOG2
`endif 

`ifdef AXI_W_S5_NMV_P1_LOG2
  `undef AXI_W_S5_NMV_P1_LOG2
`endif 

`ifdef AXI_AR_S6_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AR_S6_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AR_S6_HAS_SHRD_DDCTD_LNK
  `undef AXI_AR_S6_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AR_S6_NMV
  `undef AXI_AR_S6_NMV
`endif 

`ifdef AXI_AR_S6_NMV_LOG2
  `undef AXI_AR_S6_NMV_LOG2
`endif 

`ifdef AXI_AR_S6_NMV_P1_LOG2
  `undef AXI_AR_S6_NMV_P1_LOG2
`endif 

`ifdef AXI_AW_S6_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AW_S6_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AW_S6_HAS_SHRD_DDCTD_LNK
  `undef AXI_AW_S6_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AW_S6_NMV
  `undef AXI_AW_S6_NMV
`endif 

`ifdef AXI_AW_S6_NMV_LOG2
  `undef AXI_AW_S6_NMV_LOG2
`endif 

`ifdef AXI_AW_S6_NMV_P1_LOG2
  `undef AXI_AW_S6_NMV_P1_LOG2
`endif 

`ifdef AXI_W_S6_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_W_S6_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_W_S6_HAS_SHRD_DDCTD_LNK
  `undef AXI_W_S6_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_W_S6_NMV
  `undef AXI_W_S6_NMV
`endif 

`ifdef AXI_W_S6_NMV_LOG2
  `undef AXI_W_S6_NMV_LOG2
`endif 

`ifdef AXI_W_S6_NMV_P1_LOG2
  `undef AXI_W_S6_NMV_P1_LOG2
`endif 

`ifdef AXI_AR_S7_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AR_S7_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AR_S7_HAS_SHRD_DDCTD_LNK
  `undef AXI_AR_S7_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AR_S7_NMV
  `undef AXI_AR_S7_NMV
`endif 

`ifdef AXI_AR_S7_NMV_LOG2
  `undef AXI_AR_S7_NMV_LOG2
`endif 

`ifdef AXI_AR_S7_NMV_P1_LOG2
  `undef AXI_AR_S7_NMV_P1_LOG2
`endif 

`ifdef AXI_AW_S7_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AW_S7_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AW_S7_HAS_SHRD_DDCTD_LNK
  `undef AXI_AW_S7_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AW_S7_NMV
  `undef AXI_AW_S7_NMV
`endif 

`ifdef AXI_AW_S7_NMV_LOG2
  `undef AXI_AW_S7_NMV_LOG2
`endif 

`ifdef AXI_AW_S7_NMV_P1_LOG2
  `undef AXI_AW_S7_NMV_P1_LOG2
`endif 

`ifdef AXI_W_S7_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_W_S7_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_W_S7_HAS_SHRD_DDCTD_LNK
  `undef AXI_W_S7_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_W_S7_NMV
  `undef AXI_W_S7_NMV
`endif 

`ifdef AXI_W_S7_NMV_LOG2
  `undef AXI_W_S7_NMV_LOG2
`endif 

`ifdef AXI_W_S7_NMV_P1_LOG2
  `undef AXI_W_S7_NMV_P1_LOG2
`endif 

`ifdef AXI_AR_S8_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AR_S8_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AR_S8_HAS_SHRD_DDCTD_LNK
  `undef AXI_AR_S8_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AR_S8_NMV
  `undef AXI_AR_S8_NMV
`endif 

`ifdef AXI_AR_S8_NMV_LOG2
  `undef AXI_AR_S8_NMV_LOG2
`endif 

`ifdef AXI_AR_S8_NMV_P1_LOG2
  `undef AXI_AR_S8_NMV_P1_LOG2
`endif 

`ifdef AXI_AW_S8_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AW_S8_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AW_S8_HAS_SHRD_DDCTD_LNK
  `undef AXI_AW_S8_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AW_S8_NMV
  `undef AXI_AW_S8_NMV
`endif 

`ifdef AXI_AW_S8_NMV_LOG2
  `undef AXI_AW_S8_NMV_LOG2
`endif 

`ifdef AXI_AW_S8_NMV_P1_LOG2
  `undef AXI_AW_S8_NMV_P1_LOG2
`endif 

`ifdef AXI_W_S8_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_W_S8_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_W_S8_HAS_SHRD_DDCTD_LNK
  `undef AXI_W_S8_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_W_S8_NMV
  `undef AXI_W_S8_NMV
`endif 

`ifdef AXI_W_S8_NMV_LOG2
  `undef AXI_W_S8_NMV_LOG2
`endif 

`ifdef AXI_W_S8_NMV_P1_LOG2
  `undef AXI_W_S8_NMV_P1_LOG2
`endif 

`ifdef AXI_AR_S9_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AR_S9_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AR_S9_HAS_SHRD_DDCTD_LNK
  `undef AXI_AR_S9_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AR_S9_NMV
  `undef AXI_AR_S9_NMV
`endif 

`ifdef AXI_AR_S9_NMV_LOG2
  `undef AXI_AR_S9_NMV_LOG2
`endif 

`ifdef AXI_AR_S9_NMV_P1_LOG2
  `undef AXI_AR_S9_NMV_P1_LOG2
`endif 

`ifdef AXI_AW_S9_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AW_S9_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AW_S9_HAS_SHRD_DDCTD_LNK
  `undef AXI_AW_S9_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AW_S9_NMV
  `undef AXI_AW_S9_NMV
`endif 

`ifdef AXI_AW_S9_NMV_LOG2
  `undef AXI_AW_S9_NMV_LOG2
`endif 

`ifdef AXI_AW_S9_NMV_P1_LOG2
  `undef AXI_AW_S9_NMV_P1_LOG2
`endif 

`ifdef AXI_W_S9_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_W_S9_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_W_S9_HAS_SHRD_DDCTD_LNK
  `undef AXI_W_S9_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_W_S9_NMV
  `undef AXI_W_S9_NMV
`endif 

`ifdef AXI_W_S9_NMV_LOG2
  `undef AXI_W_S9_NMV_LOG2
`endif 

`ifdef AXI_W_S9_NMV_P1_LOG2
  `undef AXI_W_S9_NMV_P1_LOG2
`endif 

`ifdef AXI_AR_S10_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AR_S10_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AR_S10_HAS_SHRD_DDCTD_LNK
  `undef AXI_AR_S10_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AR_S10_NMV
  `undef AXI_AR_S10_NMV
`endif 

`ifdef AXI_AR_S10_NMV_LOG2
  `undef AXI_AR_S10_NMV_LOG2
`endif 

`ifdef AXI_AR_S10_NMV_P1_LOG2
  `undef AXI_AR_S10_NMV_P1_LOG2
`endif 

`ifdef AXI_AW_S10_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AW_S10_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AW_S10_HAS_SHRD_DDCTD_LNK
  `undef AXI_AW_S10_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AW_S10_NMV
  `undef AXI_AW_S10_NMV
`endif 

`ifdef AXI_AW_S10_NMV_LOG2
  `undef AXI_AW_S10_NMV_LOG2
`endif 

`ifdef AXI_AW_S10_NMV_P1_LOG2
  `undef AXI_AW_S10_NMV_P1_LOG2
`endif 

`ifdef AXI_W_S10_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_W_S10_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_W_S10_HAS_SHRD_DDCTD_LNK
  `undef AXI_W_S10_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_W_S10_NMV
  `undef AXI_W_S10_NMV
`endif 

`ifdef AXI_W_S10_NMV_LOG2
  `undef AXI_W_S10_NMV_LOG2
`endif 

`ifdef AXI_W_S10_NMV_P1_LOG2
  `undef AXI_W_S10_NMV_P1_LOG2
`endif 

`ifdef AXI_AR_S11_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AR_S11_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AR_S11_HAS_SHRD_DDCTD_LNK
  `undef AXI_AR_S11_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AR_S11_NMV
  `undef AXI_AR_S11_NMV
`endif 

`ifdef AXI_AR_S11_NMV_LOG2
  `undef AXI_AR_S11_NMV_LOG2
`endif 

`ifdef AXI_AR_S11_NMV_P1_LOG2
  `undef AXI_AR_S11_NMV_P1_LOG2
`endif 

`ifdef AXI_AW_S11_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AW_S11_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AW_S11_HAS_SHRD_DDCTD_LNK
  `undef AXI_AW_S11_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AW_S11_NMV
  `undef AXI_AW_S11_NMV
`endif 

`ifdef AXI_AW_S11_NMV_LOG2
  `undef AXI_AW_S11_NMV_LOG2
`endif 

`ifdef AXI_AW_S11_NMV_P1_LOG2
  `undef AXI_AW_S11_NMV_P1_LOG2
`endif 

`ifdef AXI_W_S11_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_W_S11_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_W_S11_HAS_SHRD_DDCTD_LNK
  `undef AXI_W_S11_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_W_S11_NMV
  `undef AXI_W_S11_NMV
`endif 

`ifdef AXI_W_S11_NMV_LOG2
  `undef AXI_W_S11_NMV_LOG2
`endif 

`ifdef AXI_W_S11_NMV_P1_LOG2
  `undef AXI_W_S11_NMV_P1_LOG2
`endif 

`ifdef AXI_AR_S12_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AR_S12_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AR_S12_HAS_SHRD_DDCTD_LNK
  `undef AXI_AR_S12_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AR_S12_NMV
  `undef AXI_AR_S12_NMV
`endif 

`ifdef AXI_AR_S12_NMV_LOG2
  `undef AXI_AR_S12_NMV_LOG2
`endif 

`ifdef AXI_AR_S12_NMV_P1_LOG2
  `undef AXI_AR_S12_NMV_P1_LOG2
`endif 

`ifdef AXI_AW_S12_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AW_S12_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AW_S12_HAS_SHRD_DDCTD_LNK
  `undef AXI_AW_S12_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AW_S12_NMV
  `undef AXI_AW_S12_NMV
`endif 

`ifdef AXI_AW_S12_NMV_LOG2
  `undef AXI_AW_S12_NMV_LOG2
`endif 

`ifdef AXI_AW_S12_NMV_P1_LOG2
  `undef AXI_AW_S12_NMV_P1_LOG2
`endif 

`ifdef AXI_W_S12_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_W_S12_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_W_S12_HAS_SHRD_DDCTD_LNK
  `undef AXI_W_S12_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_W_S12_NMV
  `undef AXI_W_S12_NMV
`endif 

`ifdef AXI_W_S12_NMV_LOG2
  `undef AXI_W_S12_NMV_LOG2
`endif 

`ifdef AXI_W_S12_NMV_P1_LOG2
  `undef AXI_W_S12_NMV_P1_LOG2
`endif 

`ifdef AXI_AR_S13_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AR_S13_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AR_S13_HAS_SHRD_DDCTD_LNK
  `undef AXI_AR_S13_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AR_S13_NMV
  `undef AXI_AR_S13_NMV
`endif 

`ifdef AXI_AR_S13_NMV_LOG2
  `undef AXI_AR_S13_NMV_LOG2
`endif 

`ifdef AXI_AR_S13_NMV_P1_LOG2
  `undef AXI_AR_S13_NMV_P1_LOG2
`endif 

`ifdef AXI_AW_S13_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AW_S13_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AW_S13_HAS_SHRD_DDCTD_LNK
  `undef AXI_AW_S13_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AW_S13_NMV
  `undef AXI_AW_S13_NMV
`endif 

`ifdef AXI_AW_S13_NMV_LOG2
  `undef AXI_AW_S13_NMV_LOG2
`endif 

`ifdef AXI_AW_S13_NMV_P1_LOG2
  `undef AXI_AW_S13_NMV_P1_LOG2
`endif 

`ifdef AXI_W_S13_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_W_S13_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_W_S13_HAS_SHRD_DDCTD_LNK
  `undef AXI_W_S13_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_W_S13_NMV
  `undef AXI_W_S13_NMV
`endif 

`ifdef AXI_W_S13_NMV_LOG2
  `undef AXI_W_S13_NMV_LOG2
`endif 

`ifdef AXI_W_S13_NMV_P1_LOG2
  `undef AXI_W_S13_NMV_P1_LOG2
`endif 

`ifdef AXI_AR_S14_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AR_S14_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AR_S14_HAS_SHRD_DDCTD_LNK
  `undef AXI_AR_S14_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AR_S14_NMV
  `undef AXI_AR_S14_NMV
`endif 

`ifdef AXI_AR_S14_NMV_LOG2
  `undef AXI_AR_S14_NMV_LOG2
`endif 

`ifdef AXI_AR_S14_NMV_P1_LOG2
  `undef AXI_AR_S14_NMV_P1_LOG2
`endif 

`ifdef AXI_AW_S14_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AW_S14_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AW_S14_HAS_SHRD_DDCTD_LNK
  `undef AXI_AW_S14_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AW_S14_NMV
  `undef AXI_AW_S14_NMV
`endif 

`ifdef AXI_AW_S14_NMV_LOG2
  `undef AXI_AW_S14_NMV_LOG2
`endif 

`ifdef AXI_AW_S14_NMV_P1_LOG2
  `undef AXI_AW_S14_NMV_P1_LOG2
`endif 

`ifdef AXI_W_S14_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_W_S14_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_W_S14_HAS_SHRD_DDCTD_LNK
  `undef AXI_W_S14_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_W_S14_NMV
  `undef AXI_W_S14_NMV
`endif 

`ifdef AXI_W_S14_NMV_LOG2
  `undef AXI_W_S14_NMV_LOG2
`endif 

`ifdef AXI_W_S14_NMV_P1_LOG2
  `undef AXI_W_S14_NMV_P1_LOG2
`endif 

`ifdef AXI_AR_S15_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AR_S15_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AR_S15_HAS_SHRD_DDCTD_LNK
  `undef AXI_AR_S15_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AR_S15_NMV
  `undef AXI_AR_S15_NMV
`endif 

`ifdef AXI_AR_S15_NMV_LOG2
  `undef AXI_AR_S15_NMV_LOG2
`endif 

`ifdef AXI_AR_S15_NMV_P1_LOG2
  `undef AXI_AR_S15_NMV_P1_LOG2
`endif 

`ifdef AXI_AW_S15_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AW_S15_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AW_S15_HAS_SHRD_DDCTD_LNK
  `undef AXI_AW_S15_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AW_S15_NMV
  `undef AXI_AW_S15_NMV
`endif 

`ifdef AXI_AW_S15_NMV_LOG2
  `undef AXI_AW_S15_NMV_LOG2
`endif 

`ifdef AXI_AW_S15_NMV_P1_LOG2
  `undef AXI_AW_S15_NMV_P1_LOG2
`endif 

`ifdef AXI_W_S15_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_W_S15_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_W_S15_HAS_SHRD_DDCTD_LNK
  `undef AXI_W_S15_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_W_S15_NMV
  `undef AXI_W_S15_NMV
`endif 

`ifdef AXI_W_S15_NMV_LOG2
  `undef AXI_W_S15_NMV_LOG2
`endif 

`ifdef AXI_W_S15_NMV_P1_LOG2
  `undef AXI_W_S15_NMV_P1_LOG2
`endif 

`ifdef AXI_AR_S16_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AR_S16_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AR_S16_HAS_SHRD_DDCTD_LNK
  `undef AXI_AR_S16_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AR_S16_NMV
  `undef AXI_AR_S16_NMV
`endif 

`ifdef AXI_AR_S16_NMV_LOG2
  `undef AXI_AR_S16_NMV_LOG2
`endif 

`ifdef AXI_AR_S16_NMV_P1_LOG2
  `undef AXI_AR_S16_NMV_P1_LOG2
`endif 

`ifdef AXI_AW_S16_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_AW_S16_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_AW_S16_HAS_SHRD_DDCTD_LNK
  `undef AXI_AW_S16_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_AW_S16_NMV
  `undef AXI_AW_S16_NMV
`endif 

`ifdef AXI_AW_S16_NMV_LOG2
  `undef AXI_AW_S16_NMV_LOG2
`endif 

`ifdef AXI_AW_S16_NMV_P1_LOG2
  `undef AXI_AW_S16_NMV_P1_LOG2
`endif 

`ifdef AXI_W_S16_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_W_S16_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_W_S16_HAS_SHRD_DDCTD_LNK
  `undef AXI_W_S16_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_W_S16_NMV
  `undef AXI_W_S16_NMV
`endif 

`ifdef AXI_W_S16_NMV_LOG2
  `undef AXI_W_S16_NMV_LOG2
`endif 

`ifdef AXI_W_S16_NMV_P1_LOG2
  `undef AXI_W_S16_NMV_P1_LOG2
`endif 

`ifdef AXI_R_M1_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_R_M1_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_R_M1_HAS_SHRD_DDCTD_LNK
  `undef AXI_R_M1_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_R_M1_NSV
  `undef AXI_R_M1_NSV
`endif 

`ifdef AXI_R_M1_NSV_LOG2
  `undef AXI_R_M1_NSV_LOG2
`endif 

`ifdef AXI_R_M1_NSV_P1_LOG2
  `undef AXI_R_M1_NSV_P1_LOG2
`endif 

`ifdef AXI_B_M1_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_B_M1_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_B_M1_HAS_SHRD_DDCTD_LNK
  `undef AXI_B_M1_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_B_M1_NSV
  `undef AXI_B_M1_NSV
`endif 

`ifdef AXI_B_M1_NSV_LOG2
  `undef AXI_B_M1_NSV_LOG2
`endif 

`ifdef AXI_B_M1_NSV_P1_LOG2
  `undef AXI_B_M1_NSV_P1_LOG2
`endif 

`ifdef AXI_R_M2_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_R_M2_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_R_M2_HAS_SHRD_DDCTD_LNK
  `undef AXI_R_M2_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_R_M2_NSV
  `undef AXI_R_M2_NSV
`endif 

`ifdef AXI_R_M2_NSV_LOG2
  `undef AXI_R_M2_NSV_LOG2
`endif 

`ifdef AXI_R_M2_NSV_P1_LOG2
  `undef AXI_R_M2_NSV_P1_LOG2
`endif 

`ifdef AXI_B_M2_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_B_M2_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_B_M2_HAS_SHRD_DDCTD_LNK
  `undef AXI_B_M2_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_B_M2_NSV
  `undef AXI_B_M2_NSV
`endif 

`ifdef AXI_B_M2_NSV_LOG2
  `undef AXI_B_M2_NSV_LOG2
`endif 

`ifdef AXI_B_M2_NSV_P1_LOG2
  `undef AXI_B_M2_NSV_P1_LOG2
`endif 

`ifdef AXI_R_M3_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_R_M3_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_R_M3_HAS_SHRD_DDCTD_LNK
  `undef AXI_R_M3_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_R_M3_NSV
  `undef AXI_R_M3_NSV
`endif 

`ifdef AXI_R_M3_NSV_LOG2
  `undef AXI_R_M3_NSV_LOG2
`endif 

`ifdef AXI_R_M3_NSV_P1_LOG2
  `undef AXI_R_M3_NSV_P1_LOG2
`endif 

`ifdef AXI_B_M3_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_B_M3_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_B_M3_HAS_SHRD_DDCTD_LNK
  `undef AXI_B_M3_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_B_M3_NSV
  `undef AXI_B_M3_NSV
`endif 

`ifdef AXI_B_M3_NSV_LOG2
  `undef AXI_B_M3_NSV_LOG2
`endif 

`ifdef AXI_B_M3_NSV_P1_LOG2
  `undef AXI_B_M3_NSV_P1_LOG2
`endif 

`ifdef AXI_R_M4_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_R_M4_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_R_M4_HAS_SHRD_DDCTD_LNK
  `undef AXI_R_M4_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_R_M4_NSV
  `undef AXI_R_M4_NSV
`endif 

`ifdef AXI_R_M4_NSV_LOG2
  `undef AXI_R_M4_NSV_LOG2
`endif 

`ifdef AXI_R_M4_NSV_P1_LOG2
  `undef AXI_R_M4_NSV_P1_LOG2
`endif 

`ifdef AXI_B_M4_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_B_M4_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_B_M4_HAS_SHRD_DDCTD_LNK
  `undef AXI_B_M4_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_B_M4_NSV
  `undef AXI_B_M4_NSV
`endif 

`ifdef AXI_B_M4_NSV_LOG2
  `undef AXI_B_M4_NSV_LOG2
`endif 

`ifdef AXI_B_M4_NSV_P1_LOG2
  `undef AXI_B_M4_NSV_P1_LOG2
`endif 

`ifdef AXI_R_M5_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_R_M5_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_R_M5_HAS_SHRD_DDCTD_LNK
  `undef AXI_R_M5_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_R_M5_NSV
  `undef AXI_R_M5_NSV
`endif 

`ifdef AXI_R_M5_NSV_LOG2
  `undef AXI_R_M5_NSV_LOG2
`endif 

`ifdef AXI_R_M5_NSV_P1_LOG2
  `undef AXI_R_M5_NSV_P1_LOG2
`endif 

`ifdef AXI_B_M5_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_B_M5_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_B_M5_HAS_SHRD_DDCTD_LNK
  `undef AXI_B_M5_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_B_M5_NSV
  `undef AXI_B_M5_NSV
`endif 

`ifdef AXI_B_M5_NSV_LOG2
  `undef AXI_B_M5_NSV_LOG2
`endif 

`ifdef AXI_B_M5_NSV_P1_LOG2
  `undef AXI_B_M5_NSV_P1_LOG2
`endif 

`ifdef AXI_R_M6_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_R_M6_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_R_M6_HAS_SHRD_DDCTD_LNK
  `undef AXI_R_M6_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_R_M6_NSV
  `undef AXI_R_M6_NSV
`endif 

`ifdef AXI_R_M6_NSV_LOG2
  `undef AXI_R_M6_NSV_LOG2
`endif 

`ifdef AXI_R_M6_NSV_P1_LOG2
  `undef AXI_R_M6_NSV_P1_LOG2
`endif 

`ifdef AXI_B_M6_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_B_M6_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_B_M6_HAS_SHRD_DDCTD_LNK
  `undef AXI_B_M6_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_B_M6_NSV
  `undef AXI_B_M6_NSV
`endif 

`ifdef AXI_B_M6_NSV_LOG2
  `undef AXI_B_M6_NSV_LOG2
`endif 

`ifdef AXI_B_M6_NSV_P1_LOG2
  `undef AXI_B_M6_NSV_P1_LOG2
`endif 

`ifdef AXI_R_M7_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_R_M7_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_R_M7_HAS_SHRD_DDCTD_LNK
  `undef AXI_R_M7_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_R_M7_NSV
  `undef AXI_R_M7_NSV
`endif 

`ifdef AXI_R_M7_NSV_LOG2
  `undef AXI_R_M7_NSV_LOG2
`endif 

`ifdef AXI_R_M7_NSV_P1_LOG2
  `undef AXI_R_M7_NSV_P1_LOG2
`endif 

`ifdef AXI_B_M7_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_B_M7_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_B_M7_HAS_SHRD_DDCTD_LNK
  `undef AXI_B_M7_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_B_M7_NSV
  `undef AXI_B_M7_NSV
`endif 

`ifdef AXI_B_M7_NSV_LOG2
  `undef AXI_B_M7_NSV_LOG2
`endif 

`ifdef AXI_B_M7_NSV_P1_LOG2
  `undef AXI_B_M7_NSV_P1_LOG2
`endif 

`ifdef AXI_R_M8_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_R_M8_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_R_M8_HAS_SHRD_DDCTD_LNK
  `undef AXI_R_M8_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_R_M8_NSV
  `undef AXI_R_M8_NSV
`endif 

`ifdef AXI_R_M8_NSV_LOG2
  `undef AXI_R_M8_NSV_LOG2
`endif 

`ifdef AXI_R_M8_NSV_P1_LOG2
  `undef AXI_R_M8_NSV_P1_LOG2
`endif 

`ifdef AXI_B_M8_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_B_M8_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_B_M8_HAS_SHRD_DDCTD_LNK
  `undef AXI_B_M8_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_B_M8_NSV
  `undef AXI_B_M8_NSV
`endif 

`ifdef AXI_B_M8_NSV_LOG2
  `undef AXI_B_M8_NSV_LOG2
`endif 

`ifdef AXI_B_M8_NSV_P1_LOG2
  `undef AXI_B_M8_NSV_P1_LOG2
`endif 

`ifdef AXI_R_M9_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_R_M9_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_R_M9_HAS_SHRD_DDCTD_LNK
  `undef AXI_R_M9_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_R_M9_NSV
  `undef AXI_R_M9_NSV
`endif 

`ifdef AXI_R_M9_NSV_LOG2
  `undef AXI_R_M9_NSV_LOG2
`endif 

`ifdef AXI_R_M9_NSV_P1_LOG2
  `undef AXI_R_M9_NSV_P1_LOG2
`endif 

`ifdef AXI_B_M9_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_B_M9_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_B_M9_HAS_SHRD_DDCTD_LNK
  `undef AXI_B_M9_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_B_M9_NSV
  `undef AXI_B_M9_NSV
`endif 

`ifdef AXI_B_M9_NSV_LOG2
  `undef AXI_B_M9_NSV_LOG2
`endif 

`ifdef AXI_B_M9_NSV_P1_LOG2
  `undef AXI_B_M9_NSV_P1_LOG2
`endif 

`ifdef AXI_R_M10_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_R_M10_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_R_M10_HAS_SHRD_DDCTD_LNK
  `undef AXI_R_M10_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_R_M10_NSV
  `undef AXI_R_M10_NSV
`endif 

`ifdef AXI_R_M10_NSV_LOG2
  `undef AXI_R_M10_NSV_LOG2
`endif 

`ifdef AXI_R_M10_NSV_P1_LOG2
  `undef AXI_R_M10_NSV_P1_LOG2
`endif 

`ifdef AXI_B_M10_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_B_M10_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_B_M10_HAS_SHRD_DDCTD_LNK
  `undef AXI_B_M10_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_B_M10_NSV
  `undef AXI_B_M10_NSV
`endif 

`ifdef AXI_B_M10_NSV_LOG2
  `undef AXI_B_M10_NSV_LOG2
`endif 

`ifdef AXI_B_M10_NSV_P1_LOG2
  `undef AXI_B_M10_NSV_P1_LOG2
`endif 

`ifdef AXI_R_M11_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_R_M11_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_R_M11_HAS_SHRD_DDCTD_LNK
  `undef AXI_R_M11_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_R_M11_NSV
  `undef AXI_R_M11_NSV
`endif 

`ifdef AXI_R_M11_NSV_LOG2
  `undef AXI_R_M11_NSV_LOG2
`endif 

`ifdef AXI_R_M11_NSV_P1_LOG2
  `undef AXI_R_M11_NSV_P1_LOG2
`endif 

`ifdef AXI_B_M11_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_B_M11_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_B_M11_HAS_SHRD_DDCTD_LNK
  `undef AXI_B_M11_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_B_M11_NSV
  `undef AXI_B_M11_NSV
`endif 

`ifdef AXI_B_M11_NSV_LOG2
  `undef AXI_B_M11_NSV_LOG2
`endif 

`ifdef AXI_B_M11_NSV_P1_LOG2
  `undef AXI_B_M11_NSV_P1_LOG2
`endif 

`ifdef AXI_R_M12_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_R_M12_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_R_M12_HAS_SHRD_DDCTD_LNK
  `undef AXI_R_M12_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_R_M12_NSV
  `undef AXI_R_M12_NSV
`endif 

`ifdef AXI_R_M12_NSV_LOG2
  `undef AXI_R_M12_NSV_LOG2
`endif 

`ifdef AXI_R_M12_NSV_P1_LOG2
  `undef AXI_R_M12_NSV_P1_LOG2
`endif 

`ifdef AXI_B_M12_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_B_M12_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_B_M12_HAS_SHRD_DDCTD_LNK
  `undef AXI_B_M12_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_B_M12_NSV
  `undef AXI_B_M12_NSV
`endif 

`ifdef AXI_B_M12_NSV_LOG2
  `undef AXI_B_M12_NSV_LOG2
`endif 

`ifdef AXI_B_M12_NSV_P1_LOG2
  `undef AXI_B_M12_NSV_P1_LOG2
`endif 

`ifdef AXI_R_M13_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_R_M13_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_R_M13_HAS_SHRD_DDCTD_LNK
  `undef AXI_R_M13_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_R_M13_NSV
  `undef AXI_R_M13_NSV
`endif 

`ifdef AXI_R_M13_NSV_LOG2
  `undef AXI_R_M13_NSV_LOG2
`endif 

`ifdef AXI_R_M13_NSV_P1_LOG2
  `undef AXI_R_M13_NSV_P1_LOG2
`endif 

`ifdef AXI_B_M13_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_B_M13_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_B_M13_HAS_SHRD_DDCTD_LNK
  `undef AXI_B_M13_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_B_M13_NSV
  `undef AXI_B_M13_NSV
`endif 

`ifdef AXI_B_M13_NSV_LOG2
  `undef AXI_B_M13_NSV_LOG2
`endif 

`ifdef AXI_B_M13_NSV_P1_LOG2
  `undef AXI_B_M13_NSV_P1_LOG2
`endif 

`ifdef AXI_R_M14_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_R_M14_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_R_M14_HAS_SHRD_DDCTD_LNK
  `undef AXI_R_M14_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_R_M14_NSV
  `undef AXI_R_M14_NSV
`endif 

`ifdef AXI_R_M14_NSV_LOG2
  `undef AXI_R_M14_NSV_LOG2
`endif 

`ifdef AXI_R_M14_NSV_P1_LOG2
  `undef AXI_R_M14_NSV_P1_LOG2
`endif 

`ifdef AXI_B_M14_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_B_M14_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_B_M14_HAS_SHRD_DDCTD_LNK
  `undef AXI_B_M14_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_B_M14_NSV
  `undef AXI_B_M14_NSV
`endif 

`ifdef AXI_B_M14_NSV_LOG2
  `undef AXI_B_M14_NSV_LOG2
`endif 

`ifdef AXI_B_M14_NSV_P1_LOG2
  `undef AXI_B_M14_NSV_P1_LOG2
`endif 

`ifdef AXI_R_M15_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_R_M15_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_R_M15_HAS_SHRD_DDCTD_LNK
  `undef AXI_R_M15_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_R_M15_NSV
  `undef AXI_R_M15_NSV
`endif 

`ifdef AXI_R_M15_NSV_LOG2
  `undef AXI_R_M15_NSV_LOG2
`endif 

`ifdef AXI_R_M15_NSV_P1_LOG2
  `undef AXI_R_M15_NSV_P1_LOG2
`endif 

`ifdef AXI_B_M15_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_B_M15_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_B_M15_HAS_SHRD_DDCTD_LNK
  `undef AXI_B_M15_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_B_M15_NSV
  `undef AXI_B_M15_NSV
`endif 

`ifdef AXI_B_M15_NSV_LOG2
  `undef AXI_B_M15_NSV_LOG2
`endif 

`ifdef AXI_B_M15_NSV_P1_LOG2
  `undef AXI_B_M15_NSV_P1_LOG2
`endif 

`ifdef AXI_R_M16_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_R_M16_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_R_M16_HAS_SHRD_DDCTD_LNK
  `undef AXI_R_M16_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_R_M16_NSV
  `undef AXI_R_M16_NSV
`endif 

`ifdef AXI_R_M16_NSV_LOG2
  `undef AXI_R_M16_NSV_LOG2
`endif 

`ifdef AXI_R_M16_NSV_P1_LOG2
  `undef AXI_R_M16_NSV_P1_LOG2
`endif 

`ifdef AXI_B_M16_HAS_SHRD_DDCTD_LNK_VAL
  `undef AXI_B_M16_HAS_SHRD_DDCTD_LNK_VAL
`endif 

`ifdef AXI_B_M16_HAS_SHRD_DDCTD_LNK
  `undef AXI_B_M16_HAS_SHRD_DDCTD_LNK
`endif 

`ifdef AXI_B_M16_NSV
  `undef AXI_B_M16_NSV
`endif 

`ifdef AXI_B_M16_NSV_LOG2
  `undef AXI_B_M16_NSV_LOG2
`endif 

`ifdef AXI_B_M16_NSV_P1_LOG2
  `undef AXI_B_M16_NSV_P1_LOG2
`endif 

`ifdef AXI_M1_ON_AR_SHARED_VAL
  `undef AXI_M1_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_M2_ON_AR_SHARED_VAL
  `undef AXI_M2_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_M3_ON_AR_SHARED_VAL
  `undef AXI_M3_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_M4_ON_AR_SHARED_VAL
  `undef AXI_M4_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_M5_ON_AR_SHARED_VAL
  `undef AXI_M5_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_M6_ON_AR_SHARED_VAL
  `undef AXI_M6_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_M7_ON_AR_SHARED_VAL
  `undef AXI_M7_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_M8_ON_AR_SHARED_VAL
  `undef AXI_M8_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_M9_ON_AR_SHARED_VAL
  `undef AXI_M9_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_M10_ON_AR_SHARED_VAL
  `undef AXI_M10_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_M11_ON_AR_SHARED_VAL
  `undef AXI_M11_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_M12_ON_AR_SHARED_VAL
  `undef AXI_M12_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_M13_ON_AR_SHARED_VAL
  `undef AXI_M13_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_M14_ON_AR_SHARED_VAL
  `undef AXI_M14_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_M15_ON_AR_SHARED_VAL
  `undef AXI_M15_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_M16_ON_AR_SHARED_VAL
  `undef AXI_M16_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_S0_ON_AR_SHARED_VAL
  `undef AXI_S0_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_S0_ON_AR_SHARED_ONLY
  `undef AXI_S0_ON_AR_SHARED_ONLY
`endif 

`ifdef AXI_S0_ON_AR_SHARED_ONLY_VAL
  `undef AXI_S0_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S1_ON_AR_SHARED_VAL
  `undef AXI_S1_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_S1_ON_AR_SHARED_ONLY
  `undef AXI_S1_ON_AR_SHARED_ONLY
`endif 

`ifdef AXI_S1_ON_AR_SHARED_ONLY_VAL
  `undef AXI_S1_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S2_ON_AR_SHARED_VAL
  `undef AXI_S2_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_S2_ON_AR_SHARED_ONLY
  `undef AXI_S2_ON_AR_SHARED_ONLY
`endif 

`ifdef AXI_S2_ON_AR_SHARED_ONLY_VAL
  `undef AXI_S2_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S3_ON_AR_SHARED_VAL
  `undef AXI_S3_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_S3_ON_AR_SHARED_ONLY
  `undef AXI_S3_ON_AR_SHARED_ONLY
`endif 

`ifdef AXI_S3_ON_AR_SHARED_ONLY_VAL
  `undef AXI_S3_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S4_ON_AR_SHARED_VAL
  `undef AXI_S4_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_S4_ON_AR_SHARED_ONLY
  `undef AXI_S4_ON_AR_SHARED_ONLY
`endif 

`ifdef AXI_S4_ON_AR_SHARED_ONLY_VAL
  `undef AXI_S4_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S5_ON_AR_SHARED_VAL
  `undef AXI_S5_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_S5_ON_AR_SHARED_ONLY
  `undef AXI_S5_ON_AR_SHARED_ONLY
`endif 

`ifdef AXI_S5_ON_AR_SHARED_ONLY_VAL
  `undef AXI_S5_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S6_ON_AR_SHARED_VAL
  `undef AXI_S6_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_S6_ON_AR_SHARED_ONLY
  `undef AXI_S6_ON_AR_SHARED_ONLY
`endif 

`ifdef AXI_S6_ON_AR_SHARED_ONLY_VAL
  `undef AXI_S6_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S7_ON_AR_SHARED_VAL
  `undef AXI_S7_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_S7_ON_AR_SHARED_ONLY
  `undef AXI_S7_ON_AR_SHARED_ONLY
`endif 

`ifdef AXI_S7_ON_AR_SHARED_ONLY_VAL
  `undef AXI_S7_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S8_ON_AR_SHARED_VAL
  `undef AXI_S8_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_S8_ON_AR_SHARED_ONLY
  `undef AXI_S8_ON_AR_SHARED_ONLY
`endif 

`ifdef AXI_S8_ON_AR_SHARED_ONLY_VAL
  `undef AXI_S8_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S9_ON_AR_SHARED_VAL
  `undef AXI_S9_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_S9_ON_AR_SHARED_ONLY
  `undef AXI_S9_ON_AR_SHARED_ONLY
`endif 

`ifdef AXI_S9_ON_AR_SHARED_ONLY_VAL
  `undef AXI_S9_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S10_ON_AR_SHARED_VAL
  `undef AXI_S10_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_S10_ON_AR_SHARED_ONLY
  `undef AXI_S10_ON_AR_SHARED_ONLY
`endif 

`ifdef AXI_S10_ON_AR_SHARED_ONLY_VAL
  `undef AXI_S10_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S11_ON_AR_SHARED_VAL
  `undef AXI_S11_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_S11_ON_AR_SHARED_ONLY
  `undef AXI_S11_ON_AR_SHARED_ONLY
`endif 

`ifdef AXI_S11_ON_AR_SHARED_ONLY_VAL
  `undef AXI_S11_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S12_ON_AR_SHARED_VAL
  `undef AXI_S12_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_S12_ON_AR_SHARED_ONLY
  `undef AXI_S12_ON_AR_SHARED_ONLY
`endif 

`ifdef AXI_S12_ON_AR_SHARED_ONLY_VAL
  `undef AXI_S12_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S13_ON_AR_SHARED_VAL
  `undef AXI_S13_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_S13_ON_AR_SHARED_ONLY
  `undef AXI_S13_ON_AR_SHARED_ONLY
`endif 

`ifdef AXI_S13_ON_AR_SHARED_ONLY_VAL
  `undef AXI_S13_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S14_ON_AR_SHARED_VAL
  `undef AXI_S14_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_S14_ON_AR_SHARED_ONLY
  `undef AXI_S14_ON_AR_SHARED_ONLY
`endif 

`ifdef AXI_S14_ON_AR_SHARED_ONLY_VAL
  `undef AXI_S14_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S15_ON_AR_SHARED_VAL
  `undef AXI_S15_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_S15_ON_AR_SHARED_ONLY
  `undef AXI_S15_ON_AR_SHARED_ONLY
`endif 

`ifdef AXI_S15_ON_AR_SHARED_ONLY_VAL
  `undef AXI_S15_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S16_ON_AR_SHARED_VAL
  `undef AXI_S16_ON_AR_SHARED_VAL
`endif 

`ifdef AXI_S16_ON_AR_SHARED_ONLY
  `undef AXI_S16_ON_AR_SHARED_ONLY
`endif 

`ifdef AXI_S16_ON_AR_SHARED_ONLY_VAL
  `undef AXI_S16_ON_AR_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M1_ON_AW_SHARED_VAL
  `undef AXI_M1_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_M2_ON_AW_SHARED_VAL
  `undef AXI_M2_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_M3_ON_AW_SHARED_VAL
  `undef AXI_M3_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_M4_ON_AW_SHARED_VAL
  `undef AXI_M4_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_M5_ON_AW_SHARED_VAL
  `undef AXI_M5_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_M6_ON_AW_SHARED_VAL
  `undef AXI_M6_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_M7_ON_AW_SHARED_VAL
  `undef AXI_M7_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_M8_ON_AW_SHARED_VAL
  `undef AXI_M8_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_M9_ON_AW_SHARED_VAL
  `undef AXI_M9_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_M10_ON_AW_SHARED_VAL
  `undef AXI_M10_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_M11_ON_AW_SHARED_VAL
  `undef AXI_M11_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_M12_ON_AW_SHARED_VAL
  `undef AXI_M12_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_M13_ON_AW_SHARED_VAL
  `undef AXI_M13_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_M14_ON_AW_SHARED_VAL
  `undef AXI_M14_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_M15_ON_AW_SHARED_VAL
  `undef AXI_M15_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_M16_ON_AW_SHARED_VAL
  `undef AXI_M16_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_S0_ON_AW_SHARED_VAL
  `undef AXI_S0_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_S0_ON_AW_SHARED_ONLY
  `undef AXI_S0_ON_AW_SHARED_ONLY
`endif 

`ifdef AXI_S0_ON_AW_SHARED_ONLY_VAL
  `undef AXI_S0_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S1_ON_AW_SHARED_VAL
  `undef AXI_S1_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_S1_ON_AW_SHARED_ONLY
  `undef AXI_S1_ON_AW_SHARED_ONLY
`endif 

`ifdef AXI_S1_ON_AW_SHARED_ONLY_VAL
  `undef AXI_S1_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S2_ON_AW_SHARED_VAL
  `undef AXI_S2_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_S2_ON_AW_SHARED_ONLY
  `undef AXI_S2_ON_AW_SHARED_ONLY
`endif 

`ifdef AXI_S2_ON_AW_SHARED_ONLY_VAL
  `undef AXI_S2_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S3_ON_AW_SHARED_VAL
  `undef AXI_S3_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_S3_ON_AW_SHARED_ONLY
  `undef AXI_S3_ON_AW_SHARED_ONLY
`endif 

`ifdef AXI_S3_ON_AW_SHARED_ONLY_VAL
  `undef AXI_S3_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S4_ON_AW_SHARED_VAL
  `undef AXI_S4_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_S4_ON_AW_SHARED_ONLY
  `undef AXI_S4_ON_AW_SHARED_ONLY
`endif 

`ifdef AXI_S4_ON_AW_SHARED_ONLY_VAL
  `undef AXI_S4_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S5_ON_AW_SHARED_VAL
  `undef AXI_S5_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_S5_ON_AW_SHARED_ONLY
  `undef AXI_S5_ON_AW_SHARED_ONLY
`endif 

`ifdef AXI_S5_ON_AW_SHARED_ONLY_VAL
  `undef AXI_S5_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S6_ON_AW_SHARED_VAL
  `undef AXI_S6_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_S6_ON_AW_SHARED_ONLY
  `undef AXI_S6_ON_AW_SHARED_ONLY
`endif 

`ifdef AXI_S6_ON_AW_SHARED_ONLY_VAL
  `undef AXI_S6_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S7_ON_AW_SHARED_VAL
  `undef AXI_S7_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_S7_ON_AW_SHARED_ONLY
  `undef AXI_S7_ON_AW_SHARED_ONLY
`endif 

`ifdef AXI_S7_ON_AW_SHARED_ONLY_VAL
  `undef AXI_S7_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S8_ON_AW_SHARED_VAL
  `undef AXI_S8_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_S8_ON_AW_SHARED_ONLY
  `undef AXI_S8_ON_AW_SHARED_ONLY
`endif 

`ifdef AXI_S8_ON_AW_SHARED_ONLY_VAL
  `undef AXI_S8_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S9_ON_AW_SHARED_VAL
  `undef AXI_S9_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_S9_ON_AW_SHARED_ONLY
  `undef AXI_S9_ON_AW_SHARED_ONLY
`endif 

`ifdef AXI_S9_ON_AW_SHARED_ONLY_VAL
  `undef AXI_S9_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S10_ON_AW_SHARED_VAL
  `undef AXI_S10_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_S10_ON_AW_SHARED_ONLY
  `undef AXI_S10_ON_AW_SHARED_ONLY
`endif 

`ifdef AXI_S10_ON_AW_SHARED_ONLY_VAL
  `undef AXI_S10_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S11_ON_AW_SHARED_VAL
  `undef AXI_S11_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_S11_ON_AW_SHARED_ONLY
  `undef AXI_S11_ON_AW_SHARED_ONLY
`endif 

`ifdef AXI_S11_ON_AW_SHARED_ONLY_VAL
  `undef AXI_S11_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S12_ON_AW_SHARED_VAL
  `undef AXI_S12_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_S12_ON_AW_SHARED_ONLY
  `undef AXI_S12_ON_AW_SHARED_ONLY
`endif 

`ifdef AXI_S12_ON_AW_SHARED_ONLY_VAL
  `undef AXI_S12_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S13_ON_AW_SHARED_VAL
  `undef AXI_S13_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_S13_ON_AW_SHARED_ONLY
  `undef AXI_S13_ON_AW_SHARED_ONLY
`endif 

`ifdef AXI_S13_ON_AW_SHARED_ONLY_VAL
  `undef AXI_S13_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S14_ON_AW_SHARED_VAL
  `undef AXI_S14_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_S14_ON_AW_SHARED_ONLY
  `undef AXI_S14_ON_AW_SHARED_ONLY
`endif 

`ifdef AXI_S14_ON_AW_SHARED_ONLY_VAL
  `undef AXI_S14_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S15_ON_AW_SHARED_VAL
  `undef AXI_S15_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_S15_ON_AW_SHARED_ONLY
  `undef AXI_S15_ON_AW_SHARED_ONLY
`endif 

`ifdef AXI_S15_ON_AW_SHARED_ONLY_VAL
  `undef AXI_S15_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S16_ON_AW_SHARED_VAL
  `undef AXI_S16_ON_AW_SHARED_VAL
`endif 

`ifdef AXI_S16_ON_AW_SHARED_ONLY
  `undef AXI_S16_ON_AW_SHARED_ONLY
`endif 

`ifdef AXI_S16_ON_AW_SHARED_ONLY_VAL
  `undef AXI_S16_ON_AW_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M1_ON_W_SHARED_VAL
  `undef AXI_M1_ON_W_SHARED_VAL
`endif 

`ifdef AXI_M2_ON_W_SHARED_VAL
  `undef AXI_M2_ON_W_SHARED_VAL
`endif 

`ifdef AXI_M3_ON_W_SHARED_VAL
  `undef AXI_M3_ON_W_SHARED_VAL
`endif 

`ifdef AXI_M4_ON_W_SHARED_VAL
  `undef AXI_M4_ON_W_SHARED_VAL
`endif 

`ifdef AXI_M5_ON_W_SHARED_VAL
  `undef AXI_M5_ON_W_SHARED_VAL
`endif 

`ifdef AXI_M6_ON_W_SHARED_VAL
  `undef AXI_M6_ON_W_SHARED_VAL
`endif 

`ifdef AXI_M7_ON_W_SHARED_VAL
  `undef AXI_M7_ON_W_SHARED_VAL
`endif 

`ifdef AXI_M8_ON_W_SHARED_VAL
  `undef AXI_M8_ON_W_SHARED_VAL
`endif 

`ifdef AXI_M9_ON_W_SHARED_VAL
  `undef AXI_M9_ON_W_SHARED_VAL
`endif 

`ifdef AXI_M10_ON_W_SHARED_VAL
  `undef AXI_M10_ON_W_SHARED_VAL
`endif 

`ifdef AXI_M11_ON_W_SHARED_VAL
  `undef AXI_M11_ON_W_SHARED_VAL
`endif 

`ifdef AXI_M12_ON_W_SHARED_VAL
  `undef AXI_M12_ON_W_SHARED_VAL
`endif 

`ifdef AXI_M13_ON_W_SHARED_VAL
  `undef AXI_M13_ON_W_SHARED_VAL
`endif 

`ifdef AXI_M14_ON_W_SHARED_VAL
  `undef AXI_M14_ON_W_SHARED_VAL
`endif 

`ifdef AXI_M15_ON_W_SHARED_VAL
  `undef AXI_M15_ON_W_SHARED_VAL
`endif 

`ifdef AXI_M16_ON_W_SHARED_VAL
  `undef AXI_M16_ON_W_SHARED_VAL
`endif 

`ifdef AXI_S0_ON_W_SHARED_VAL
  `undef AXI_S0_ON_W_SHARED_VAL
`endif 

`ifdef AXI_S0_ON_W_SHARED_ONLY
  `undef AXI_S0_ON_W_SHARED_ONLY
`endif 

`ifdef AXI_S0_ON_W_SHARED_ONLY_VAL
  `undef AXI_S0_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S1_ON_W_SHARED_VAL
  `undef AXI_S1_ON_W_SHARED_VAL
`endif 

`ifdef AXI_S1_ON_W_SHARED_ONLY
  `undef AXI_S1_ON_W_SHARED_ONLY
`endif 

`ifdef AXI_S1_ON_W_SHARED_ONLY_VAL
  `undef AXI_S1_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S2_ON_W_SHARED_VAL
  `undef AXI_S2_ON_W_SHARED_VAL
`endif 

`ifdef AXI_S2_ON_W_SHARED_ONLY
  `undef AXI_S2_ON_W_SHARED_ONLY
`endif 

`ifdef AXI_S2_ON_W_SHARED_ONLY_VAL
  `undef AXI_S2_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S3_ON_W_SHARED_VAL
  `undef AXI_S3_ON_W_SHARED_VAL
`endif 

`ifdef AXI_S3_ON_W_SHARED_ONLY
  `undef AXI_S3_ON_W_SHARED_ONLY
`endif 

`ifdef AXI_S3_ON_W_SHARED_ONLY_VAL
  `undef AXI_S3_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S4_ON_W_SHARED_VAL
  `undef AXI_S4_ON_W_SHARED_VAL
`endif 

`ifdef AXI_S4_ON_W_SHARED_ONLY
  `undef AXI_S4_ON_W_SHARED_ONLY
`endif 

`ifdef AXI_S4_ON_W_SHARED_ONLY_VAL
  `undef AXI_S4_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S5_ON_W_SHARED_VAL
  `undef AXI_S5_ON_W_SHARED_VAL
`endif 

`ifdef AXI_S5_ON_W_SHARED_ONLY
  `undef AXI_S5_ON_W_SHARED_ONLY
`endif 

`ifdef AXI_S5_ON_W_SHARED_ONLY_VAL
  `undef AXI_S5_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S6_ON_W_SHARED_VAL
  `undef AXI_S6_ON_W_SHARED_VAL
`endif 

`ifdef AXI_S6_ON_W_SHARED_ONLY
  `undef AXI_S6_ON_W_SHARED_ONLY
`endif 

`ifdef AXI_S6_ON_W_SHARED_ONLY_VAL
  `undef AXI_S6_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S7_ON_W_SHARED_VAL
  `undef AXI_S7_ON_W_SHARED_VAL
`endif 

`ifdef AXI_S7_ON_W_SHARED_ONLY
  `undef AXI_S7_ON_W_SHARED_ONLY
`endif 

`ifdef AXI_S7_ON_W_SHARED_ONLY_VAL
  `undef AXI_S7_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S8_ON_W_SHARED_VAL
  `undef AXI_S8_ON_W_SHARED_VAL
`endif 

`ifdef AXI_S8_ON_W_SHARED_ONLY
  `undef AXI_S8_ON_W_SHARED_ONLY
`endif 

`ifdef AXI_S8_ON_W_SHARED_ONLY_VAL
  `undef AXI_S8_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S9_ON_W_SHARED_VAL
  `undef AXI_S9_ON_W_SHARED_VAL
`endif 

`ifdef AXI_S9_ON_W_SHARED_ONLY
  `undef AXI_S9_ON_W_SHARED_ONLY
`endif 

`ifdef AXI_S9_ON_W_SHARED_ONLY_VAL
  `undef AXI_S9_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S10_ON_W_SHARED_VAL
  `undef AXI_S10_ON_W_SHARED_VAL
`endif 

`ifdef AXI_S10_ON_W_SHARED_ONLY
  `undef AXI_S10_ON_W_SHARED_ONLY
`endif 

`ifdef AXI_S10_ON_W_SHARED_ONLY_VAL
  `undef AXI_S10_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S11_ON_W_SHARED_VAL
  `undef AXI_S11_ON_W_SHARED_VAL
`endif 

`ifdef AXI_S11_ON_W_SHARED_ONLY
  `undef AXI_S11_ON_W_SHARED_ONLY
`endif 

`ifdef AXI_S11_ON_W_SHARED_ONLY_VAL
  `undef AXI_S11_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S12_ON_W_SHARED_VAL
  `undef AXI_S12_ON_W_SHARED_VAL
`endif 

`ifdef AXI_S12_ON_W_SHARED_ONLY
  `undef AXI_S12_ON_W_SHARED_ONLY
`endif 

`ifdef AXI_S12_ON_W_SHARED_ONLY_VAL
  `undef AXI_S12_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S13_ON_W_SHARED_VAL
  `undef AXI_S13_ON_W_SHARED_VAL
`endif 

`ifdef AXI_S13_ON_W_SHARED_ONLY
  `undef AXI_S13_ON_W_SHARED_ONLY
`endif 

`ifdef AXI_S13_ON_W_SHARED_ONLY_VAL
  `undef AXI_S13_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S14_ON_W_SHARED_VAL
  `undef AXI_S14_ON_W_SHARED_VAL
`endif 

`ifdef AXI_S14_ON_W_SHARED_ONLY
  `undef AXI_S14_ON_W_SHARED_ONLY
`endif 

`ifdef AXI_S14_ON_W_SHARED_ONLY_VAL
  `undef AXI_S14_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S15_ON_W_SHARED_VAL
  `undef AXI_S15_ON_W_SHARED_VAL
`endif 

`ifdef AXI_S15_ON_W_SHARED_ONLY
  `undef AXI_S15_ON_W_SHARED_ONLY
`endif 

`ifdef AXI_S15_ON_W_SHARED_ONLY_VAL
  `undef AXI_S15_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S16_ON_W_SHARED_VAL
  `undef AXI_S16_ON_W_SHARED_VAL
`endif 

`ifdef AXI_S16_ON_W_SHARED_ONLY
  `undef AXI_S16_ON_W_SHARED_ONLY
`endif 

`ifdef AXI_S16_ON_W_SHARED_ONLY_VAL
  `undef AXI_S16_ON_W_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S0_ON_R_SHARED_VAL
  `undef AXI_S0_ON_R_SHARED_VAL
`endif 

`ifdef AXI_S1_ON_R_SHARED_VAL
  `undef AXI_S1_ON_R_SHARED_VAL
`endif 

`ifdef AXI_S2_ON_R_SHARED_VAL
  `undef AXI_S2_ON_R_SHARED_VAL
`endif 

`ifdef AXI_S3_ON_R_SHARED_VAL
  `undef AXI_S3_ON_R_SHARED_VAL
`endif 

`ifdef AXI_S4_ON_R_SHARED_VAL
  `undef AXI_S4_ON_R_SHARED_VAL
`endif 

`ifdef AXI_S5_ON_R_SHARED_VAL
  `undef AXI_S5_ON_R_SHARED_VAL
`endif 

`ifdef AXI_S6_ON_R_SHARED_VAL
  `undef AXI_S6_ON_R_SHARED_VAL
`endif 

`ifdef AXI_S7_ON_R_SHARED_VAL
  `undef AXI_S7_ON_R_SHARED_VAL
`endif 

`ifdef AXI_S8_ON_R_SHARED_VAL
  `undef AXI_S8_ON_R_SHARED_VAL
`endif 

`ifdef AXI_S9_ON_R_SHARED_VAL
  `undef AXI_S9_ON_R_SHARED_VAL
`endif 

`ifdef AXI_S10_ON_R_SHARED_VAL
  `undef AXI_S10_ON_R_SHARED_VAL
`endif 

`ifdef AXI_S11_ON_R_SHARED_VAL
  `undef AXI_S11_ON_R_SHARED_VAL
`endif 

`ifdef AXI_S12_ON_R_SHARED_VAL
  `undef AXI_S12_ON_R_SHARED_VAL
`endif 

`ifdef AXI_S13_ON_R_SHARED_VAL
  `undef AXI_S13_ON_R_SHARED_VAL
`endif 

`ifdef AXI_S14_ON_R_SHARED_VAL
  `undef AXI_S14_ON_R_SHARED_VAL
`endif 

`ifdef AXI_S15_ON_R_SHARED_VAL
  `undef AXI_S15_ON_R_SHARED_VAL
`endif 

`ifdef AXI_S16_ON_R_SHARED_VAL
  `undef AXI_S16_ON_R_SHARED_VAL
`endif 

`ifdef AXI_M1_ON_R_SHARED_VAL
  `undef AXI_M1_ON_R_SHARED_VAL
`endif 

`ifdef AXI_M1_ON_R_SHARED_ONLY
  `undef AXI_M1_ON_R_SHARED_ONLY
`endif 

`ifdef AXI_M1_ON_R_SHARED_ONLY_VAL
  `undef AXI_M1_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M2_ON_R_SHARED_VAL
  `undef AXI_M2_ON_R_SHARED_VAL
`endif 

`ifdef AXI_M2_ON_R_SHARED_ONLY
  `undef AXI_M2_ON_R_SHARED_ONLY
`endif 

`ifdef AXI_M2_ON_R_SHARED_ONLY_VAL
  `undef AXI_M2_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M3_ON_R_SHARED_VAL
  `undef AXI_M3_ON_R_SHARED_VAL
`endif 

`ifdef AXI_M3_ON_R_SHARED_ONLY
  `undef AXI_M3_ON_R_SHARED_ONLY
`endif 

`ifdef AXI_M3_ON_R_SHARED_ONLY_VAL
  `undef AXI_M3_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M4_ON_R_SHARED_VAL
  `undef AXI_M4_ON_R_SHARED_VAL
`endif 

`ifdef AXI_M4_ON_R_SHARED_ONLY
  `undef AXI_M4_ON_R_SHARED_ONLY
`endif 

`ifdef AXI_M4_ON_R_SHARED_ONLY_VAL
  `undef AXI_M4_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M5_ON_R_SHARED_VAL
  `undef AXI_M5_ON_R_SHARED_VAL
`endif 

`ifdef AXI_M5_ON_R_SHARED_ONLY
  `undef AXI_M5_ON_R_SHARED_ONLY
`endif 

`ifdef AXI_M5_ON_R_SHARED_ONLY_VAL
  `undef AXI_M5_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M6_ON_R_SHARED_VAL
  `undef AXI_M6_ON_R_SHARED_VAL
`endif 

`ifdef AXI_M6_ON_R_SHARED_ONLY
  `undef AXI_M6_ON_R_SHARED_ONLY
`endif 

`ifdef AXI_M6_ON_R_SHARED_ONLY_VAL
  `undef AXI_M6_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M7_ON_R_SHARED_VAL
  `undef AXI_M7_ON_R_SHARED_VAL
`endif 

`ifdef AXI_M7_ON_R_SHARED_ONLY
  `undef AXI_M7_ON_R_SHARED_ONLY
`endif 

`ifdef AXI_M7_ON_R_SHARED_ONLY_VAL
  `undef AXI_M7_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M8_ON_R_SHARED_VAL
  `undef AXI_M8_ON_R_SHARED_VAL
`endif 

`ifdef AXI_M8_ON_R_SHARED_ONLY
  `undef AXI_M8_ON_R_SHARED_ONLY
`endif 

`ifdef AXI_M8_ON_R_SHARED_ONLY_VAL
  `undef AXI_M8_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M9_ON_R_SHARED_VAL
  `undef AXI_M9_ON_R_SHARED_VAL
`endif 

`ifdef AXI_M9_ON_R_SHARED_ONLY
  `undef AXI_M9_ON_R_SHARED_ONLY
`endif 

`ifdef AXI_M9_ON_R_SHARED_ONLY_VAL
  `undef AXI_M9_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M10_ON_R_SHARED_VAL
  `undef AXI_M10_ON_R_SHARED_VAL
`endif 

`ifdef AXI_M10_ON_R_SHARED_ONLY
  `undef AXI_M10_ON_R_SHARED_ONLY
`endif 

`ifdef AXI_M10_ON_R_SHARED_ONLY_VAL
  `undef AXI_M10_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M11_ON_R_SHARED_VAL
  `undef AXI_M11_ON_R_SHARED_VAL
`endif 

`ifdef AXI_M11_ON_R_SHARED_ONLY
  `undef AXI_M11_ON_R_SHARED_ONLY
`endif 

`ifdef AXI_M11_ON_R_SHARED_ONLY_VAL
  `undef AXI_M11_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M12_ON_R_SHARED_VAL
  `undef AXI_M12_ON_R_SHARED_VAL
`endif 

`ifdef AXI_M12_ON_R_SHARED_ONLY
  `undef AXI_M12_ON_R_SHARED_ONLY
`endif 

`ifdef AXI_M12_ON_R_SHARED_ONLY_VAL
  `undef AXI_M12_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M13_ON_R_SHARED_VAL
  `undef AXI_M13_ON_R_SHARED_VAL
`endif 

`ifdef AXI_M13_ON_R_SHARED_ONLY
  `undef AXI_M13_ON_R_SHARED_ONLY
`endif 

`ifdef AXI_M13_ON_R_SHARED_ONLY_VAL
  `undef AXI_M13_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M14_ON_R_SHARED_VAL
  `undef AXI_M14_ON_R_SHARED_VAL
`endif 

`ifdef AXI_M14_ON_R_SHARED_ONLY
  `undef AXI_M14_ON_R_SHARED_ONLY
`endif 

`ifdef AXI_M14_ON_R_SHARED_ONLY_VAL
  `undef AXI_M14_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M15_ON_R_SHARED_VAL
  `undef AXI_M15_ON_R_SHARED_VAL
`endif 

`ifdef AXI_M15_ON_R_SHARED_ONLY
  `undef AXI_M15_ON_R_SHARED_ONLY
`endif 

`ifdef AXI_M15_ON_R_SHARED_ONLY_VAL
  `undef AXI_M15_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M16_ON_R_SHARED_VAL
  `undef AXI_M16_ON_R_SHARED_VAL
`endif 

`ifdef AXI_M16_ON_R_SHARED_ONLY
  `undef AXI_M16_ON_R_SHARED_ONLY
`endif 

`ifdef AXI_M16_ON_R_SHARED_ONLY_VAL
  `undef AXI_M16_ON_R_SHARED_ONLY_VAL
`endif 

`ifdef AXI_S0_ON_B_SHARED_VAL
  `undef AXI_S0_ON_B_SHARED_VAL
`endif 

`ifdef AXI_S1_ON_B_SHARED_VAL
  `undef AXI_S1_ON_B_SHARED_VAL
`endif 

`ifdef AXI_S2_ON_B_SHARED_VAL
  `undef AXI_S2_ON_B_SHARED_VAL
`endif 

`ifdef AXI_S3_ON_B_SHARED_VAL
  `undef AXI_S3_ON_B_SHARED_VAL
`endif 

`ifdef AXI_S4_ON_B_SHARED_VAL
  `undef AXI_S4_ON_B_SHARED_VAL
`endif 

`ifdef AXI_S5_ON_B_SHARED_VAL
  `undef AXI_S5_ON_B_SHARED_VAL
`endif 

`ifdef AXI_S6_ON_B_SHARED_VAL
  `undef AXI_S6_ON_B_SHARED_VAL
`endif 

`ifdef AXI_S7_ON_B_SHARED_VAL
  `undef AXI_S7_ON_B_SHARED_VAL
`endif 

`ifdef AXI_S8_ON_B_SHARED_VAL
  `undef AXI_S8_ON_B_SHARED_VAL
`endif 

`ifdef AXI_S9_ON_B_SHARED_VAL
  `undef AXI_S9_ON_B_SHARED_VAL
`endif 

`ifdef AXI_S10_ON_B_SHARED_VAL
  `undef AXI_S10_ON_B_SHARED_VAL
`endif 

`ifdef AXI_S11_ON_B_SHARED_VAL
  `undef AXI_S11_ON_B_SHARED_VAL
`endif 

`ifdef AXI_S12_ON_B_SHARED_VAL
  `undef AXI_S12_ON_B_SHARED_VAL
`endif 

`ifdef AXI_S13_ON_B_SHARED_VAL
  `undef AXI_S13_ON_B_SHARED_VAL
`endif 

`ifdef AXI_S14_ON_B_SHARED_VAL
  `undef AXI_S14_ON_B_SHARED_VAL
`endif 

`ifdef AXI_S15_ON_B_SHARED_VAL
  `undef AXI_S15_ON_B_SHARED_VAL
`endif 

`ifdef AXI_S16_ON_B_SHARED_VAL
  `undef AXI_S16_ON_B_SHARED_VAL
`endif 

`ifdef AXI_M1_ON_B_SHARED_VAL
  `undef AXI_M1_ON_B_SHARED_VAL
`endif 

`ifdef AXI_M1_ON_B_SHARED_ONLY
  `undef AXI_M1_ON_B_SHARED_ONLY
`endif 

`ifdef AXI_M1_ON_B_SHARED_ONLY_VAL
  `undef AXI_M1_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M2_ON_B_SHARED_VAL
  `undef AXI_M2_ON_B_SHARED_VAL
`endif 

`ifdef AXI_M2_ON_B_SHARED_ONLY
  `undef AXI_M2_ON_B_SHARED_ONLY
`endif 

`ifdef AXI_M2_ON_B_SHARED_ONLY_VAL
  `undef AXI_M2_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M3_ON_B_SHARED_VAL
  `undef AXI_M3_ON_B_SHARED_VAL
`endif 

`ifdef AXI_M3_ON_B_SHARED_ONLY
  `undef AXI_M3_ON_B_SHARED_ONLY
`endif 

`ifdef AXI_M3_ON_B_SHARED_ONLY_VAL
  `undef AXI_M3_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M4_ON_B_SHARED_VAL
  `undef AXI_M4_ON_B_SHARED_VAL
`endif 

`ifdef AXI_M4_ON_B_SHARED_ONLY
  `undef AXI_M4_ON_B_SHARED_ONLY
`endif 

`ifdef AXI_M4_ON_B_SHARED_ONLY_VAL
  `undef AXI_M4_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M5_ON_B_SHARED_VAL
  `undef AXI_M5_ON_B_SHARED_VAL
`endif 

`ifdef AXI_M5_ON_B_SHARED_ONLY
  `undef AXI_M5_ON_B_SHARED_ONLY
`endif 

`ifdef AXI_M5_ON_B_SHARED_ONLY_VAL
  `undef AXI_M5_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M6_ON_B_SHARED_VAL
  `undef AXI_M6_ON_B_SHARED_VAL
`endif 

`ifdef AXI_M6_ON_B_SHARED_ONLY
  `undef AXI_M6_ON_B_SHARED_ONLY
`endif 

`ifdef AXI_M6_ON_B_SHARED_ONLY_VAL
  `undef AXI_M6_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M7_ON_B_SHARED_VAL
  `undef AXI_M7_ON_B_SHARED_VAL
`endif 

`ifdef AXI_M7_ON_B_SHARED_ONLY
  `undef AXI_M7_ON_B_SHARED_ONLY
`endif 

`ifdef AXI_M7_ON_B_SHARED_ONLY_VAL
  `undef AXI_M7_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M8_ON_B_SHARED_VAL
  `undef AXI_M8_ON_B_SHARED_VAL
`endif 

`ifdef AXI_M8_ON_B_SHARED_ONLY
  `undef AXI_M8_ON_B_SHARED_ONLY
`endif 

`ifdef AXI_M8_ON_B_SHARED_ONLY_VAL
  `undef AXI_M8_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M9_ON_B_SHARED_VAL
  `undef AXI_M9_ON_B_SHARED_VAL
`endif 

`ifdef AXI_M9_ON_B_SHARED_ONLY
  `undef AXI_M9_ON_B_SHARED_ONLY
`endif 

`ifdef AXI_M9_ON_B_SHARED_ONLY_VAL
  `undef AXI_M9_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M10_ON_B_SHARED_VAL
  `undef AXI_M10_ON_B_SHARED_VAL
`endif 

`ifdef AXI_M10_ON_B_SHARED_ONLY
  `undef AXI_M10_ON_B_SHARED_ONLY
`endif 

`ifdef AXI_M10_ON_B_SHARED_ONLY_VAL
  `undef AXI_M10_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M11_ON_B_SHARED_VAL
  `undef AXI_M11_ON_B_SHARED_VAL
`endif 

`ifdef AXI_M11_ON_B_SHARED_ONLY
  `undef AXI_M11_ON_B_SHARED_ONLY
`endif 

`ifdef AXI_M11_ON_B_SHARED_ONLY_VAL
  `undef AXI_M11_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M12_ON_B_SHARED_VAL
  `undef AXI_M12_ON_B_SHARED_VAL
`endif 

`ifdef AXI_M12_ON_B_SHARED_ONLY
  `undef AXI_M12_ON_B_SHARED_ONLY
`endif 

`ifdef AXI_M12_ON_B_SHARED_ONLY_VAL
  `undef AXI_M12_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M13_ON_B_SHARED_VAL
  `undef AXI_M13_ON_B_SHARED_VAL
`endif 

`ifdef AXI_M13_ON_B_SHARED_ONLY
  `undef AXI_M13_ON_B_SHARED_ONLY
`endif 

`ifdef AXI_M13_ON_B_SHARED_ONLY_VAL
  `undef AXI_M13_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M14_ON_B_SHARED_VAL
  `undef AXI_M14_ON_B_SHARED_VAL
`endif 

`ifdef AXI_M14_ON_B_SHARED_ONLY
  `undef AXI_M14_ON_B_SHARED_ONLY
`endif 

`ifdef AXI_M14_ON_B_SHARED_ONLY_VAL
  `undef AXI_M14_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M15_ON_B_SHARED_VAL
  `undef AXI_M15_ON_B_SHARED_VAL
`endif 

`ifdef AXI_M15_ON_B_SHARED_ONLY
  `undef AXI_M15_ON_B_SHARED_ONLY
`endif 

`ifdef AXI_M15_ON_B_SHARED_ONLY_VAL
  `undef AXI_M15_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef AXI_M16_ON_B_SHARED_VAL
  `undef AXI_M16_ON_B_SHARED_VAL
`endif 

`ifdef AXI_M16_ON_B_SHARED_ONLY
  `undef AXI_M16_ON_B_SHARED_ONLY
`endif 

`ifdef AXI_M16_ON_B_SHARED_ONLY_VAL
  `undef AXI_M16_ON_B_SHARED_ONLY_VAL
`endif 

`ifdef AXI_AW_SHARED_PL
  `undef AXI_AW_SHARED_PL
`endif 

`ifdef AXI_AR_SHARED_PL
  `undef AXI_AR_SHARED_PL
`endif 

`ifdef AXI_W_SHARED_PL
  `undef AXI_W_SHARED_PL
`endif 

`ifdef AXI_R_SHARED_PL
  `undef AXI_R_SHARED_PL
`endif 

`ifdef AXI_B_SHARED_PL
  `undef AXI_B_SHARED_PL
`endif 

`ifdef AXI_MCA_HLD_PRIOR
  `undef AXI_MCA_HLD_PRIOR
`endif 

`ifdef AXI_AR_MCA_NC_S0
  `undef AXI_AR_MCA_NC_S0
`endif 

`ifdef AXI_AR_MCA_EN_S0
  `undef AXI_AR_MCA_EN_S0
`endif 

`ifdef AXI_AR_MCA_NC_W_S0
  `undef AXI_AR_MCA_NC_W_S0
`endif 

`ifdef AXI_AW_MCA_NC_S0
  `undef AXI_AW_MCA_NC_S0
`endif 

`ifdef AXI_AW_MCA_EN_S0
  `undef AXI_AW_MCA_EN_S0
`endif 

`ifdef AXI_AW_MCA_NC_W_S0
  `undef AXI_AW_MCA_NC_W_S0
`endif 

`ifdef AXI_W_MCA_NC_S0
  `undef AXI_W_MCA_NC_S0
`endif 

`ifdef AXI_W_MCA_EN_S0
  `undef AXI_W_MCA_EN_S0
`endif 

`ifdef AXI_W_MCA_NC_W_S0
  `undef AXI_W_MCA_NC_W_S0
`endif 

`ifdef AXI_AR_MCA_NC_S1
  `undef AXI_AR_MCA_NC_S1
`endif 

`ifdef AXI_AR_MCA_EN_S1
  `undef AXI_AR_MCA_EN_S1
`endif 

`ifdef AXI_AR_MCA_NC_W_S1
  `undef AXI_AR_MCA_NC_W_S1
`endif 

`ifdef AXI_AW_MCA_NC_S1
  `undef AXI_AW_MCA_NC_S1
`endif 

`ifdef AXI_AW_MCA_EN_S1
  `undef AXI_AW_MCA_EN_S1
`endif 

`ifdef AXI_AW_MCA_NC_W_S1
  `undef AXI_AW_MCA_NC_W_S1
`endif 

`ifdef AXI_W_MCA_NC_S1
  `undef AXI_W_MCA_NC_S1
`endif 

`ifdef AXI_W_MCA_EN_S1
  `undef AXI_W_MCA_EN_S1
`endif 

`ifdef AXI_W_MCA_NC_W_S1
  `undef AXI_W_MCA_NC_W_S1
`endif 

`ifdef AXI_AR_MCA_NC_S2
  `undef AXI_AR_MCA_NC_S2
`endif 

`ifdef AXI_AR_MCA_EN_S2
  `undef AXI_AR_MCA_EN_S2
`endif 

`ifdef AXI_AR_MCA_NC_W_S2
  `undef AXI_AR_MCA_NC_W_S2
`endif 

`ifdef AXI_AW_MCA_NC_S2
  `undef AXI_AW_MCA_NC_S2
`endif 

`ifdef AXI_AW_MCA_EN_S2
  `undef AXI_AW_MCA_EN_S2
`endif 

`ifdef AXI_AW_MCA_NC_W_S2
  `undef AXI_AW_MCA_NC_W_S2
`endif 

`ifdef AXI_W_MCA_NC_S2
  `undef AXI_W_MCA_NC_S2
`endif 

`ifdef AXI_W_MCA_EN_S2
  `undef AXI_W_MCA_EN_S2
`endif 

`ifdef AXI_W_MCA_NC_W_S2
  `undef AXI_W_MCA_NC_W_S2
`endif 

`ifdef AXI_AR_MCA_NC_S3
  `undef AXI_AR_MCA_NC_S3
`endif 

`ifdef AXI_AR_MCA_EN_S3
  `undef AXI_AR_MCA_EN_S3
`endif 

`ifdef AXI_AR_MCA_NC_W_S3
  `undef AXI_AR_MCA_NC_W_S3
`endif 

`ifdef AXI_AW_MCA_NC_S3
  `undef AXI_AW_MCA_NC_S3
`endif 

`ifdef AXI_AW_MCA_EN_S3
  `undef AXI_AW_MCA_EN_S3
`endif 

`ifdef AXI_AW_MCA_NC_W_S3
  `undef AXI_AW_MCA_NC_W_S3
`endif 

`ifdef AXI_W_MCA_NC_S3
  `undef AXI_W_MCA_NC_S3
`endif 

`ifdef AXI_W_MCA_EN_S3
  `undef AXI_W_MCA_EN_S3
`endif 

`ifdef AXI_W_MCA_NC_W_S3
  `undef AXI_W_MCA_NC_W_S3
`endif 

`ifdef AXI_AR_MCA_NC_S4
  `undef AXI_AR_MCA_NC_S4
`endif 

`ifdef AXI_AR_MCA_EN_S4
  `undef AXI_AR_MCA_EN_S4
`endif 

`ifdef AXI_AR_MCA_NC_W_S4
  `undef AXI_AR_MCA_NC_W_S4
`endif 

`ifdef AXI_AW_MCA_NC_S4
  `undef AXI_AW_MCA_NC_S4
`endif 

`ifdef AXI_AW_MCA_EN_S4
  `undef AXI_AW_MCA_EN_S4
`endif 

`ifdef AXI_AW_MCA_NC_W_S4
  `undef AXI_AW_MCA_NC_W_S4
`endif 

`ifdef AXI_W_MCA_NC_S4
  `undef AXI_W_MCA_NC_S4
`endif 

`ifdef AXI_W_MCA_EN_S4
  `undef AXI_W_MCA_EN_S4
`endif 

`ifdef AXI_W_MCA_NC_W_S4
  `undef AXI_W_MCA_NC_W_S4
`endif 

`ifdef AXI_AR_MCA_NC_S5
  `undef AXI_AR_MCA_NC_S5
`endif 

`ifdef AXI_AR_MCA_EN_S5
  `undef AXI_AR_MCA_EN_S5
`endif 

`ifdef AXI_AR_MCA_NC_W_S5
  `undef AXI_AR_MCA_NC_W_S5
`endif 

`ifdef AXI_AW_MCA_NC_S5
  `undef AXI_AW_MCA_NC_S5
`endif 

`ifdef AXI_AW_MCA_EN_S5
  `undef AXI_AW_MCA_EN_S5
`endif 

`ifdef AXI_AW_MCA_NC_W_S5
  `undef AXI_AW_MCA_NC_W_S5
`endif 

`ifdef AXI_W_MCA_NC_S5
  `undef AXI_W_MCA_NC_S5
`endif 

`ifdef AXI_W_MCA_EN_S5
  `undef AXI_W_MCA_EN_S5
`endif 

`ifdef AXI_W_MCA_NC_W_S5
  `undef AXI_W_MCA_NC_W_S5
`endif 

`ifdef AXI_AR_MCA_NC_S6
  `undef AXI_AR_MCA_NC_S6
`endif 

`ifdef AXI_AR_MCA_EN_S6
  `undef AXI_AR_MCA_EN_S6
`endif 

`ifdef AXI_AR_MCA_NC_W_S6
  `undef AXI_AR_MCA_NC_W_S6
`endif 

`ifdef AXI_AW_MCA_NC_S6
  `undef AXI_AW_MCA_NC_S6
`endif 

`ifdef AXI_AW_MCA_EN_S6
  `undef AXI_AW_MCA_EN_S6
`endif 

`ifdef AXI_AW_MCA_NC_W_S6
  `undef AXI_AW_MCA_NC_W_S6
`endif 

`ifdef AXI_W_MCA_NC_S6
  `undef AXI_W_MCA_NC_S6
`endif 

`ifdef AXI_W_MCA_EN_S6
  `undef AXI_W_MCA_EN_S6
`endif 

`ifdef AXI_W_MCA_NC_W_S6
  `undef AXI_W_MCA_NC_W_S6
`endif 

`ifdef AXI_AR_MCA_NC_S7
  `undef AXI_AR_MCA_NC_S7
`endif 

`ifdef AXI_AR_MCA_EN_S7
  `undef AXI_AR_MCA_EN_S7
`endif 

`ifdef AXI_AR_MCA_NC_W_S7
  `undef AXI_AR_MCA_NC_W_S7
`endif 

`ifdef AXI_AW_MCA_NC_S7
  `undef AXI_AW_MCA_NC_S7
`endif 

`ifdef AXI_AW_MCA_EN_S7
  `undef AXI_AW_MCA_EN_S7
`endif 

`ifdef AXI_AW_MCA_NC_W_S7
  `undef AXI_AW_MCA_NC_W_S7
`endif 

`ifdef AXI_W_MCA_NC_S7
  `undef AXI_W_MCA_NC_S7
`endif 

`ifdef AXI_W_MCA_EN_S7
  `undef AXI_W_MCA_EN_S7
`endif 

`ifdef AXI_W_MCA_NC_W_S7
  `undef AXI_W_MCA_NC_W_S7
`endif 

`ifdef AXI_AR_MCA_NC_S8
  `undef AXI_AR_MCA_NC_S8
`endif 

`ifdef AXI_AR_MCA_EN_S8
  `undef AXI_AR_MCA_EN_S8
`endif 

`ifdef AXI_AR_MCA_NC_W_S8
  `undef AXI_AR_MCA_NC_W_S8
`endif 

`ifdef AXI_AW_MCA_NC_S8
  `undef AXI_AW_MCA_NC_S8
`endif 

`ifdef AXI_AW_MCA_EN_S8
  `undef AXI_AW_MCA_EN_S8
`endif 

`ifdef AXI_AW_MCA_NC_W_S8
  `undef AXI_AW_MCA_NC_W_S8
`endif 

`ifdef AXI_W_MCA_NC_S8
  `undef AXI_W_MCA_NC_S8
`endif 

`ifdef AXI_W_MCA_EN_S8
  `undef AXI_W_MCA_EN_S8
`endif 

`ifdef AXI_W_MCA_NC_W_S8
  `undef AXI_W_MCA_NC_W_S8
`endif 

`ifdef AXI_AR_MCA_NC_S9
  `undef AXI_AR_MCA_NC_S9
`endif 

`ifdef AXI_AR_MCA_EN_S9
  `undef AXI_AR_MCA_EN_S9
`endif 

`ifdef AXI_AR_MCA_NC_W_S9
  `undef AXI_AR_MCA_NC_W_S9
`endif 

`ifdef AXI_AW_MCA_NC_S9
  `undef AXI_AW_MCA_NC_S9
`endif 

`ifdef AXI_AW_MCA_EN_S9
  `undef AXI_AW_MCA_EN_S9
`endif 

`ifdef AXI_AW_MCA_NC_W_S9
  `undef AXI_AW_MCA_NC_W_S9
`endif 

`ifdef AXI_W_MCA_NC_S9
  `undef AXI_W_MCA_NC_S9
`endif 

`ifdef AXI_W_MCA_EN_S9
  `undef AXI_W_MCA_EN_S9
`endif 

`ifdef AXI_W_MCA_NC_W_S9
  `undef AXI_W_MCA_NC_W_S9
`endif 

`ifdef AXI_AR_MCA_NC_S10
  `undef AXI_AR_MCA_NC_S10
`endif 

`ifdef AXI_AR_MCA_EN_S10
  `undef AXI_AR_MCA_EN_S10
`endif 

`ifdef AXI_AR_MCA_NC_W_S10
  `undef AXI_AR_MCA_NC_W_S10
`endif 

`ifdef AXI_AW_MCA_NC_S10
  `undef AXI_AW_MCA_NC_S10
`endif 

`ifdef AXI_AW_MCA_EN_S10
  `undef AXI_AW_MCA_EN_S10
`endif 

`ifdef AXI_AW_MCA_NC_W_S10
  `undef AXI_AW_MCA_NC_W_S10
`endif 

`ifdef AXI_W_MCA_NC_S10
  `undef AXI_W_MCA_NC_S10
`endif 

`ifdef AXI_W_MCA_EN_S10
  `undef AXI_W_MCA_EN_S10
`endif 

`ifdef AXI_W_MCA_NC_W_S10
  `undef AXI_W_MCA_NC_W_S10
`endif 

`ifdef AXI_AR_MCA_NC_S11
  `undef AXI_AR_MCA_NC_S11
`endif 

`ifdef AXI_AR_MCA_EN_S11
  `undef AXI_AR_MCA_EN_S11
`endif 

`ifdef AXI_AR_MCA_NC_W_S11
  `undef AXI_AR_MCA_NC_W_S11
`endif 

`ifdef AXI_AW_MCA_NC_S11
  `undef AXI_AW_MCA_NC_S11
`endif 

`ifdef AXI_AW_MCA_EN_S11
  `undef AXI_AW_MCA_EN_S11
`endif 

`ifdef AXI_AW_MCA_NC_W_S11
  `undef AXI_AW_MCA_NC_W_S11
`endif 

`ifdef AXI_W_MCA_NC_S11
  `undef AXI_W_MCA_NC_S11
`endif 

`ifdef AXI_W_MCA_EN_S11
  `undef AXI_W_MCA_EN_S11
`endif 

`ifdef AXI_W_MCA_NC_W_S11
  `undef AXI_W_MCA_NC_W_S11
`endif 

`ifdef AXI_AR_MCA_NC_S12
  `undef AXI_AR_MCA_NC_S12
`endif 

`ifdef AXI_AR_MCA_EN_S12
  `undef AXI_AR_MCA_EN_S12
`endif 

`ifdef AXI_AR_MCA_NC_W_S12
  `undef AXI_AR_MCA_NC_W_S12
`endif 

`ifdef AXI_AW_MCA_NC_S12
  `undef AXI_AW_MCA_NC_S12
`endif 

`ifdef AXI_AW_MCA_EN_S12
  `undef AXI_AW_MCA_EN_S12
`endif 

`ifdef AXI_AW_MCA_NC_W_S12
  `undef AXI_AW_MCA_NC_W_S12
`endif 

`ifdef AXI_W_MCA_NC_S12
  `undef AXI_W_MCA_NC_S12
`endif 

`ifdef AXI_W_MCA_EN_S12
  `undef AXI_W_MCA_EN_S12
`endif 

`ifdef AXI_W_MCA_NC_W_S12
  `undef AXI_W_MCA_NC_W_S12
`endif 

`ifdef AXI_AR_MCA_NC_S13
  `undef AXI_AR_MCA_NC_S13
`endif 

`ifdef AXI_AR_MCA_EN_S13
  `undef AXI_AR_MCA_EN_S13
`endif 

`ifdef AXI_AR_MCA_NC_W_S13
  `undef AXI_AR_MCA_NC_W_S13
`endif 

`ifdef AXI_AW_MCA_NC_S13
  `undef AXI_AW_MCA_NC_S13
`endif 

`ifdef AXI_AW_MCA_EN_S13
  `undef AXI_AW_MCA_EN_S13
`endif 

`ifdef AXI_AW_MCA_NC_W_S13
  `undef AXI_AW_MCA_NC_W_S13
`endif 

`ifdef AXI_W_MCA_NC_S13
  `undef AXI_W_MCA_NC_S13
`endif 

`ifdef AXI_W_MCA_EN_S13
  `undef AXI_W_MCA_EN_S13
`endif 

`ifdef AXI_W_MCA_NC_W_S13
  `undef AXI_W_MCA_NC_W_S13
`endif 

`ifdef AXI_AR_MCA_NC_S14
  `undef AXI_AR_MCA_NC_S14
`endif 

`ifdef AXI_AR_MCA_EN_S14
  `undef AXI_AR_MCA_EN_S14
`endif 

`ifdef AXI_AR_MCA_NC_W_S14
  `undef AXI_AR_MCA_NC_W_S14
`endif 

`ifdef AXI_AW_MCA_NC_S14
  `undef AXI_AW_MCA_NC_S14
`endif 

`ifdef AXI_AW_MCA_EN_S14
  `undef AXI_AW_MCA_EN_S14
`endif 

`ifdef AXI_AW_MCA_NC_W_S14
  `undef AXI_AW_MCA_NC_W_S14
`endif 

`ifdef AXI_W_MCA_NC_S14
  `undef AXI_W_MCA_NC_S14
`endif 

`ifdef AXI_W_MCA_EN_S14
  `undef AXI_W_MCA_EN_S14
`endif 

`ifdef AXI_W_MCA_NC_W_S14
  `undef AXI_W_MCA_NC_W_S14
`endif 

`ifdef AXI_AR_MCA_NC_S15
  `undef AXI_AR_MCA_NC_S15
`endif 

`ifdef AXI_AR_MCA_EN_S15
  `undef AXI_AR_MCA_EN_S15
`endif 

`ifdef AXI_AR_MCA_NC_W_S15
  `undef AXI_AR_MCA_NC_W_S15
`endif 

`ifdef AXI_AW_MCA_NC_S15
  `undef AXI_AW_MCA_NC_S15
`endif 

`ifdef AXI_AW_MCA_EN_S15
  `undef AXI_AW_MCA_EN_S15
`endif 

`ifdef AXI_AW_MCA_NC_W_S15
  `undef AXI_AW_MCA_NC_W_S15
`endif 

`ifdef AXI_W_MCA_NC_S15
  `undef AXI_W_MCA_NC_S15
`endif 

`ifdef AXI_W_MCA_EN_S15
  `undef AXI_W_MCA_EN_S15
`endif 

`ifdef AXI_W_MCA_NC_W_S15
  `undef AXI_W_MCA_NC_W_S15
`endif 

`ifdef AXI_AR_MCA_NC_S16
  `undef AXI_AR_MCA_NC_S16
`endif 

`ifdef AXI_AR_MCA_EN_S16
  `undef AXI_AR_MCA_EN_S16
`endif 

`ifdef AXI_AR_MCA_NC_W_S16
  `undef AXI_AR_MCA_NC_W_S16
`endif 

`ifdef AXI_AW_MCA_NC_S16
  `undef AXI_AW_MCA_NC_S16
`endif 

`ifdef AXI_AW_MCA_EN_S16
  `undef AXI_AW_MCA_EN_S16
`endif 

`ifdef AXI_AW_MCA_NC_W_S16
  `undef AXI_AW_MCA_NC_W_S16
`endif 

`ifdef AXI_W_MCA_NC_S16
  `undef AXI_W_MCA_NC_S16
`endif 

`ifdef AXI_W_MCA_EN_S16
  `undef AXI_W_MCA_EN_S16
`endif 

`ifdef AXI_W_MCA_NC_W_S16
  `undef AXI_W_MCA_NC_W_S16
`endif 

`ifdef AXI_R_MCA_NC_M1
  `undef AXI_R_MCA_NC_M1
`endif 

`ifdef AXI_R_MCA_EN_M1
  `undef AXI_R_MCA_EN_M1
`endif 

`ifdef AXI_R_MCA_NC_W_M1
  `undef AXI_R_MCA_NC_W_M1
`endif 

`ifdef AXI_B_MCA_NC_M1
  `undef AXI_B_MCA_NC_M1
`endif 

`ifdef AXI_B_MCA_EN_M1
  `undef AXI_B_MCA_EN_M1
`endif 

`ifdef AXI_B_MCA_NC_W_M1
  `undef AXI_B_MCA_NC_W_M1
`endif 

`ifdef AXI_R_MCA_NC_M2
  `undef AXI_R_MCA_NC_M2
`endif 

`ifdef AXI_R_MCA_EN_M2
  `undef AXI_R_MCA_EN_M2
`endif 

`ifdef AXI_R_MCA_NC_W_M2
  `undef AXI_R_MCA_NC_W_M2
`endif 

`ifdef AXI_B_MCA_NC_M2
  `undef AXI_B_MCA_NC_M2
`endif 

`ifdef AXI_B_MCA_EN_M2
  `undef AXI_B_MCA_EN_M2
`endif 

`ifdef AXI_B_MCA_NC_W_M2
  `undef AXI_B_MCA_NC_W_M2
`endif 

`ifdef AXI_R_MCA_NC_M3
  `undef AXI_R_MCA_NC_M3
`endif 

`ifdef AXI_R_MCA_EN_M3
  `undef AXI_R_MCA_EN_M3
`endif 

`ifdef AXI_R_MCA_NC_W_M3
  `undef AXI_R_MCA_NC_W_M3
`endif 

`ifdef AXI_B_MCA_NC_M3
  `undef AXI_B_MCA_NC_M3
`endif 

`ifdef AXI_B_MCA_EN_M3
  `undef AXI_B_MCA_EN_M3
`endif 

`ifdef AXI_B_MCA_NC_W_M3
  `undef AXI_B_MCA_NC_W_M3
`endif 

`ifdef AXI_R_MCA_NC_M4
  `undef AXI_R_MCA_NC_M4
`endif 

`ifdef AXI_R_MCA_EN_M4
  `undef AXI_R_MCA_EN_M4
`endif 

`ifdef AXI_R_MCA_NC_W_M4
  `undef AXI_R_MCA_NC_W_M4
`endif 

`ifdef AXI_B_MCA_NC_M4
  `undef AXI_B_MCA_NC_M4
`endif 

`ifdef AXI_B_MCA_EN_M4
  `undef AXI_B_MCA_EN_M4
`endif 

`ifdef AXI_B_MCA_NC_W_M4
  `undef AXI_B_MCA_NC_W_M4
`endif 

`ifdef AXI_R_MCA_NC_M5
  `undef AXI_R_MCA_NC_M5
`endif 

`ifdef AXI_R_MCA_EN_M5
  `undef AXI_R_MCA_EN_M5
`endif 

`ifdef AXI_R_MCA_NC_W_M5
  `undef AXI_R_MCA_NC_W_M5
`endif 

`ifdef AXI_B_MCA_NC_M5
  `undef AXI_B_MCA_NC_M5
`endif 

`ifdef AXI_B_MCA_EN_M5
  `undef AXI_B_MCA_EN_M5
`endif 

`ifdef AXI_B_MCA_NC_W_M5
  `undef AXI_B_MCA_NC_W_M5
`endif 

`ifdef AXI_R_MCA_NC_M6
  `undef AXI_R_MCA_NC_M6
`endif 

`ifdef AXI_R_MCA_EN_M6
  `undef AXI_R_MCA_EN_M6
`endif 

`ifdef AXI_R_MCA_NC_W_M6
  `undef AXI_R_MCA_NC_W_M6
`endif 

`ifdef AXI_B_MCA_NC_M6
  `undef AXI_B_MCA_NC_M6
`endif 

`ifdef AXI_B_MCA_EN_M6
  `undef AXI_B_MCA_EN_M6
`endif 

`ifdef AXI_B_MCA_NC_W_M6
  `undef AXI_B_MCA_NC_W_M6
`endif 

`ifdef AXI_R_MCA_NC_M7
  `undef AXI_R_MCA_NC_M7
`endif 

`ifdef AXI_R_MCA_EN_M7
  `undef AXI_R_MCA_EN_M7
`endif 

`ifdef AXI_R_MCA_NC_W_M7
  `undef AXI_R_MCA_NC_W_M7
`endif 

`ifdef AXI_B_MCA_NC_M7
  `undef AXI_B_MCA_NC_M7
`endif 

`ifdef AXI_B_MCA_EN_M7
  `undef AXI_B_MCA_EN_M7
`endif 

`ifdef AXI_B_MCA_NC_W_M7
  `undef AXI_B_MCA_NC_W_M7
`endif 

`ifdef AXI_R_MCA_NC_M8
  `undef AXI_R_MCA_NC_M8
`endif 

`ifdef AXI_R_MCA_EN_M8
  `undef AXI_R_MCA_EN_M8
`endif 

`ifdef AXI_R_MCA_NC_W_M8
  `undef AXI_R_MCA_NC_W_M8
`endif 

`ifdef AXI_B_MCA_NC_M8
  `undef AXI_B_MCA_NC_M8
`endif 

`ifdef AXI_B_MCA_EN_M8
  `undef AXI_B_MCA_EN_M8
`endif 

`ifdef AXI_B_MCA_NC_W_M8
  `undef AXI_B_MCA_NC_W_M8
`endif 

`ifdef AXI_R_MCA_NC_M9
  `undef AXI_R_MCA_NC_M9
`endif 

`ifdef AXI_R_MCA_EN_M9
  `undef AXI_R_MCA_EN_M9
`endif 

`ifdef AXI_R_MCA_NC_W_M9
  `undef AXI_R_MCA_NC_W_M9
`endif 

`ifdef AXI_B_MCA_NC_M9
  `undef AXI_B_MCA_NC_M9
`endif 

`ifdef AXI_B_MCA_EN_M9
  `undef AXI_B_MCA_EN_M9
`endif 

`ifdef AXI_B_MCA_NC_W_M9
  `undef AXI_B_MCA_NC_W_M9
`endif 

`ifdef AXI_R_MCA_NC_M10
  `undef AXI_R_MCA_NC_M10
`endif 

`ifdef AXI_R_MCA_EN_M10
  `undef AXI_R_MCA_EN_M10
`endif 

`ifdef AXI_R_MCA_NC_W_M10
  `undef AXI_R_MCA_NC_W_M10
`endif 

`ifdef AXI_B_MCA_NC_M10
  `undef AXI_B_MCA_NC_M10
`endif 

`ifdef AXI_B_MCA_EN_M10
  `undef AXI_B_MCA_EN_M10
`endif 

`ifdef AXI_B_MCA_NC_W_M10
  `undef AXI_B_MCA_NC_W_M10
`endif 

`ifdef AXI_R_MCA_NC_M11
  `undef AXI_R_MCA_NC_M11
`endif 

`ifdef AXI_R_MCA_EN_M11
  `undef AXI_R_MCA_EN_M11
`endif 

`ifdef AXI_R_MCA_NC_W_M11
  `undef AXI_R_MCA_NC_W_M11
`endif 

`ifdef AXI_B_MCA_NC_M11
  `undef AXI_B_MCA_NC_M11
`endif 

`ifdef AXI_B_MCA_EN_M11
  `undef AXI_B_MCA_EN_M11
`endif 

`ifdef AXI_B_MCA_NC_W_M11
  `undef AXI_B_MCA_NC_W_M11
`endif 

`ifdef AXI_R_MCA_NC_M12
  `undef AXI_R_MCA_NC_M12
`endif 

`ifdef AXI_R_MCA_EN_M12
  `undef AXI_R_MCA_EN_M12
`endif 

`ifdef AXI_R_MCA_NC_W_M12
  `undef AXI_R_MCA_NC_W_M12
`endif 

`ifdef AXI_B_MCA_NC_M12
  `undef AXI_B_MCA_NC_M12
`endif 

`ifdef AXI_B_MCA_EN_M12
  `undef AXI_B_MCA_EN_M12
`endif 

`ifdef AXI_B_MCA_NC_W_M12
  `undef AXI_B_MCA_NC_W_M12
`endif 

`ifdef AXI_R_MCA_NC_M13
  `undef AXI_R_MCA_NC_M13
`endif 

`ifdef AXI_R_MCA_EN_M13
  `undef AXI_R_MCA_EN_M13
`endif 

`ifdef AXI_R_MCA_NC_W_M13
  `undef AXI_R_MCA_NC_W_M13
`endif 

`ifdef AXI_B_MCA_NC_M13
  `undef AXI_B_MCA_NC_M13
`endif 

`ifdef AXI_B_MCA_EN_M13
  `undef AXI_B_MCA_EN_M13
`endif 

`ifdef AXI_B_MCA_NC_W_M13
  `undef AXI_B_MCA_NC_W_M13
`endif 

`ifdef AXI_R_MCA_NC_M14
  `undef AXI_R_MCA_NC_M14
`endif 

`ifdef AXI_R_MCA_EN_M14
  `undef AXI_R_MCA_EN_M14
`endif 

`ifdef AXI_R_MCA_NC_W_M14
  `undef AXI_R_MCA_NC_W_M14
`endif 

`ifdef AXI_B_MCA_NC_M14
  `undef AXI_B_MCA_NC_M14
`endif 

`ifdef AXI_B_MCA_EN_M14
  `undef AXI_B_MCA_EN_M14
`endif 

`ifdef AXI_B_MCA_NC_W_M14
  `undef AXI_B_MCA_NC_W_M14
`endif 

`ifdef AXI_R_MCA_NC_M15
  `undef AXI_R_MCA_NC_M15
`endif 

`ifdef AXI_R_MCA_EN_M15
  `undef AXI_R_MCA_EN_M15
`endif 

`ifdef AXI_R_MCA_NC_W_M15
  `undef AXI_R_MCA_NC_W_M15
`endif 

`ifdef AXI_B_MCA_NC_M15
  `undef AXI_B_MCA_NC_M15
`endif 

`ifdef AXI_B_MCA_EN_M15
  `undef AXI_B_MCA_EN_M15
`endif 

`ifdef AXI_B_MCA_NC_W_M15
  `undef AXI_B_MCA_NC_W_M15
`endif 

`ifdef AXI_R_MCA_NC_M16
  `undef AXI_R_MCA_NC_M16
`endif 

`ifdef AXI_R_MCA_EN_M16
  `undef AXI_R_MCA_EN_M16
`endif 

`ifdef AXI_R_MCA_NC_W_M16
  `undef AXI_R_MCA_NC_W_M16
`endif 

`ifdef AXI_B_MCA_NC_M16
  `undef AXI_B_MCA_NC_M16
`endif 

`ifdef AXI_B_MCA_EN_M16
  `undef AXI_B_MCA_EN_M16
`endif 

`ifdef AXI_B_MCA_NC_W_M16
  `undef AXI_B_MCA_NC_W_M16
`endif 

`ifdef AXI_AR_SHARED_MCA_NC
  `undef AXI_AR_SHARED_MCA_NC
`endif 

`ifdef AXI_AR_SHARED_MCA_EN
  `undef AXI_AR_SHARED_MCA_EN
`endif 

`ifdef AXI_AR_SHARED_MCA_NC_W
  `undef AXI_AR_SHARED_MCA_NC_W
`endif 

`ifdef AXI_AW_SHARED_MCA_NC
  `undef AXI_AW_SHARED_MCA_NC
`endif 

`ifdef AXI_AW_SHARED_MCA_EN
  `undef AXI_AW_SHARED_MCA_EN
`endif 

`ifdef AXI_AW_SHARED_MCA_NC_W
  `undef AXI_AW_SHARED_MCA_NC_W
`endif 

`ifdef AXI_W_SHARED_MCA_NC
  `undef AXI_W_SHARED_MCA_NC
`endif 

`ifdef AXI_W_SHARED_MCA_EN
  `undef AXI_W_SHARED_MCA_EN
`endif 

`ifdef AXI_W_SHARED_MCA_NC_W
  `undef AXI_W_SHARED_MCA_NC_W
`endif 

`ifdef AXI_R_SHARED_MCA_NC
  `undef AXI_R_SHARED_MCA_NC
`endif 

`ifdef AXI_R_SHARED_MCA_EN
  `undef AXI_R_SHARED_MCA_EN
`endif 

`ifdef AXI_R_SHARED_MCA_NC_W
  `undef AXI_R_SHARED_MCA_NC_W
`endif 

`ifdef AXI_B_SHARED_MCA_NC
  `undef AXI_B_SHARED_MCA_NC
`endif 

`ifdef AXI_B_SHARED_MCA_EN
  `undef AXI_B_SHARED_MCA_EN
`endif 

`ifdef AXI_B_SHARED_MCA_NC_W
  `undef AXI_B_SHARED_MCA_NC_W
`endif 

`ifdef AXI_MAX_RCA_ID_M1
  `undef AXI_MAX_RCA_ID_M1
`endif 

`ifdef AXI_LOG2_MAX_RCA_ID_P1_M1
  `undef AXI_LOG2_MAX_RCA_ID_P1_M1
`endif 

`ifdef AXI_MAX_WCA_ID_M1
  `undef AXI_MAX_WCA_ID_M1
`endif 

`ifdef AXI_LOG2_MAX_WCA_ID_P1_M1
  `undef AXI_LOG2_MAX_WCA_ID_P1_M1
`endif 

`ifdef AXI_MAX_URIDA_M1
  `undef AXI_MAX_URIDA_M1
`endif 

`ifdef AXI_LOG2_MAX_URIDA_M1
  `undef AXI_LOG2_MAX_URIDA_M1
`endif 

`ifdef AXI_MAX_UWIDA_M1
  `undef AXI_MAX_UWIDA_M1
`endif 

`ifdef AXI_LOG2_MAX_UWIDA_M1
  `undef AXI_LOG2_MAX_UWIDA_M1
`endif 

`ifdef AXI_RI_LIMIT_M1
  `undef AXI_RI_LIMIT_M1
`endif 

`ifdef AXI_MAX_RCA_ID_M2
  `undef AXI_MAX_RCA_ID_M2
`endif 

`ifdef AXI_LOG2_MAX_RCA_ID_P1_M2
  `undef AXI_LOG2_MAX_RCA_ID_P1_M2
`endif 

`ifdef AXI_MAX_WCA_ID_M2
  `undef AXI_MAX_WCA_ID_M2
`endif 

`ifdef AXI_LOG2_MAX_WCA_ID_P1_M2
  `undef AXI_LOG2_MAX_WCA_ID_P1_M2
`endif 

`ifdef AXI_MAX_URIDA_M2
  `undef AXI_MAX_URIDA_M2
`endif 

`ifdef AXI_LOG2_MAX_URIDA_M2
  `undef AXI_LOG2_MAX_URIDA_M2
`endif 

`ifdef AXI_MAX_UWIDA_M2
  `undef AXI_MAX_UWIDA_M2
`endif 

`ifdef AXI_LOG2_MAX_UWIDA_M2
  `undef AXI_LOG2_MAX_UWIDA_M2
`endif 

`ifdef AXI_RI_LIMIT_M2
  `undef AXI_RI_LIMIT_M2
`endif 

`ifdef AXI_MAX_RCA_ID_M3
  `undef AXI_MAX_RCA_ID_M3
`endif 

`ifdef AXI_LOG2_MAX_RCA_ID_P1_M3
  `undef AXI_LOG2_MAX_RCA_ID_P1_M3
`endif 

`ifdef AXI_MAX_WCA_ID_M3
  `undef AXI_MAX_WCA_ID_M3
`endif 

`ifdef AXI_LOG2_MAX_WCA_ID_P1_M3
  `undef AXI_LOG2_MAX_WCA_ID_P1_M3
`endif 

`ifdef AXI_MAX_URIDA_M3
  `undef AXI_MAX_URIDA_M3
`endif 

`ifdef AXI_LOG2_MAX_URIDA_M3
  `undef AXI_LOG2_MAX_URIDA_M3
`endif 

`ifdef AXI_MAX_UWIDA_M3
  `undef AXI_MAX_UWIDA_M3
`endif 

`ifdef AXI_LOG2_MAX_UWIDA_M3
  `undef AXI_LOG2_MAX_UWIDA_M3
`endif 

`ifdef AXI_RI_LIMIT_M3
  `undef AXI_RI_LIMIT_M3
`endif 

`ifdef AXI_MAX_RCA_ID_M4
  `undef AXI_MAX_RCA_ID_M4
`endif 

`ifdef AXI_LOG2_MAX_RCA_ID_P1_M4
  `undef AXI_LOG2_MAX_RCA_ID_P1_M4
`endif 

`ifdef AXI_MAX_WCA_ID_M4
  `undef AXI_MAX_WCA_ID_M4
`endif 

`ifdef AXI_LOG2_MAX_WCA_ID_P1_M4
  `undef AXI_LOG2_MAX_WCA_ID_P1_M4
`endif 

`ifdef AXI_MAX_URIDA_M4
  `undef AXI_MAX_URIDA_M4
`endif 

`ifdef AXI_LOG2_MAX_URIDA_M4
  `undef AXI_LOG2_MAX_URIDA_M4
`endif 

`ifdef AXI_MAX_UWIDA_M4
  `undef AXI_MAX_UWIDA_M4
`endif 

`ifdef AXI_LOG2_MAX_UWIDA_M4
  `undef AXI_LOG2_MAX_UWIDA_M4
`endif 

`ifdef AXI_RI_LIMIT_M4
  `undef AXI_RI_LIMIT_M4
`endif 

`ifdef AXI_MAX_RCA_ID_M5
  `undef AXI_MAX_RCA_ID_M5
`endif 

`ifdef AXI_LOG2_MAX_RCA_ID_P1_M5
  `undef AXI_LOG2_MAX_RCA_ID_P1_M5
`endif 

`ifdef AXI_MAX_WCA_ID_M5
  `undef AXI_MAX_WCA_ID_M5
`endif 

`ifdef AXI_LOG2_MAX_WCA_ID_P1_M5
  `undef AXI_LOG2_MAX_WCA_ID_P1_M5
`endif 

`ifdef AXI_MAX_URIDA_M5
  `undef AXI_MAX_URIDA_M5
`endif 

`ifdef AXI_LOG2_MAX_URIDA_M5
  `undef AXI_LOG2_MAX_URIDA_M5
`endif 

`ifdef AXI_MAX_UWIDA_M5
  `undef AXI_MAX_UWIDA_M5
`endif 

`ifdef AXI_LOG2_MAX_UWIDA_M5
  `undef AXI_LOG2_MAX_UWIDA_M5
`endif 

`ifdef AXI_RI_LIMIT_M5
  `undef AXI_RI_LIMIT_M5
`endif 

`ifdef AXI_MAX_RCA_ID_M6
  `undef AXI_MAX_RCA_ID_M6
`endif 

`ifdef AXI_LOG2_MAX_RCA_ID_P1_M6
  `undef AXI_LOG2_MAX_RCA_ID_P1_M6
`endif 

`ifdef AXI_MAX_WCA_ID_M6
  `undef AXI_MAX_WCA_ID_M6
`endif 

`ifdef AXI_LOG2_MAX_WCA_ID_P1_M6
  `undef AXI_LOG2_MAX_WCA_ID_P1_M6
`endif 

`ifdef AXI_MAX_URIDA_M6
  `undef AXI_MAX_URIDA_M6
`endif 

`ifdef AXI_LOG2_MAX_URIDA_M6
  `undef AXI_LOG2_MAX_URIDA_M6
`endif 

`ifdef AXI_MAX_UWIDA_M6
  `undef AXI_MAX_UWIDA_M6
`endif 

`ifdef AXI_LOG2_MAX_UWIDA_M6
  `undef AXI_LOG2_MAX_UWIDA_M6
`endif 

`ifdef AXI_RI_LIMIT_M6
  `undef AXI_RI_LIMIT_M6
`endif 

`ifdef AXI_MAX_RCA_ID_M7
  `undef AXI_MAX_RCA_ID_M7
`endif 

`ifdef AXI_LOG2_MAX_RCA_ID_P1_M7
  `undef AXI_LOG2_MAX_RCA_ID_P1_M7
`endif 

`ifdef AXI_MAX_WCA_ID_M7
  `undef AXI_MAX_WCA_ID_M7
`endif 

`ifdef AXI_LOG2_MAX_WCA_ID_P1_M7
  `undef AXI_LOG2_MAX_WCA_ID_P1_M7
`endif 

`ifdef AXI_MAX_URIDA_M7
  `undef AXI_MAX_URIDA_M7
`endif 

`ifdef AXI_LOG2_MAX_URIDA_M7
  `undef AXI_LOG2_MAX_URIDA_M7
`endif 

`ifdef AXI_MAX_UWIDA_M7
  `undef AXI_MAX_UWIDA_M7
`endif 

`ifdef AXI_LOG2_MAX_UWIDA_M7
  `undef AXI_LOG2_MAX_UWIDA_M7
`endif 

`ifdef AXI_RI_LIMIT_M7
  `undef AXI_RI_LIMIT_M7
`endif 

`ifdef AXI_MAX_RCA_ID_M8
  `undef AXI_MAX_RCA_ID_M8
`endif 

`ifdef AXI_LOG2_MAX_RCA_ID_P1_M8
  `undef AXI_LOG2_MAX_RCA_ID_P1_M8
`endif 

`ifdef AXI_MAX_WCA_ID_M8
  `undef AXI_MAX_WCA_ID_M8
`endif 

`ifdef AXI_LOG2_MAX_WCA_ID_P1_M8
  `undef AXI_LOG2_MAX_WCA_ID_P1_M8
`endif 

`ifdef AXI_MAX_URIDA_M8
  `undef AXI_MAX_URIDA_M8
`endif 

`ifdef AXI_LOG2_MAX_URIDA_M8
  `undef AXI_LOG2_MAX_URIDA_M8
`endif 

`ifdef AXI_MAX_UWIDA_M8
  `undef AXI_MAX_UWIDA_M8
`endif 

`ifdef AXI_LOG2_MAX_UWIDA_M8
  `undef AXI_LOG2_MAX_UWIDA_M8
`endif 

`ifdef AXI_RI_LIMIT_M8
  `undef AXI_RI_LIMIT_M8
`endif 

`ifdef AXI_MAX_RCA_ID_M9
  `undef AXI_MAX_RCA_ID_M9
`endif 

`ifdef AXI_LOG2_MAX_RCA_ID_P1_M9
  `undef AXI_LOG2_MAX_RCA_ID_P1_M9
`endif 

`ifdef AXI_MAX_WCA_ID_M9
  `undef AXI_MAX_WCA_ID_M9
`endif 

`ifdef AXI_LOG2_MAX_WCA_ID_P1_M9
  `undef AXI_LOG2_MAX_WCA_ID_P1_M9
`endif 

`ifdef AXI_MAX_URIDA_M9
  `undef AXI_MAX_URIDA_M9
`endif 

`ifdef AXI_LOG2_MAX_URIDA_M9
  `undef AXI_LOG2_MAX_URIDA_M9
`endif 

`ifdef AXI_MAX_UWIDA_M9
  `undef AXI_MAX_UWIDA_M9
`endif 

`ifdef AXI_LOG2_MAX_UWIDA_M9
  `undef AXI_LOG2_MAX_UWIDA_M9
`endif 

`ifdef AXI_RI_LIMIT_M9
  `undef AXI_RI_LIMIT_M9
`endif 

`ifdef AXI_MAX_RCA_ID_M10
  `undef AXI_MAX_RCA_ID_M10
`endif 

`ifdef AXI_LOG2_MAX_RCA_ID_P1_M10
  `undef AXI_LOG2_MAX_RCA_ID_P1_M10
`endif 

`ifdef AXI_MAX_WCA_ID_M10
  `undef AXI_MAX_WCA_ID_M10
`endif 

`ifdef AXI_LOG2_MAX_WCA_ID_P1_M10
  `undef AXI_LOG2_MAX_WCA_ID_P1_M10
`endif 

`ifdef AXI_MAX_URIDA_M10
  `undef AXI_MAX_URIDA_M10
`endif 

`ifdef AXI_LOG2_MAX_URIDA_M10
  `undef AXI_LOG2_MAX_URIDA_M10
`endif 

`ifdef AXI_MAX_UWIDA_M10
  `undef AXI_MAX_UWIDA_M10
`endif 

`ifdef AXI_LOG2_MAX_UWIDA_M10
  `undef AXI_LOG2_MAX_UWIDA_M10
`endif 

`ifdef AXI_RI_LIMIT_M10
  `undef AXI_RI_LIMIT_M10
`endif 

`ifdef AXI_MAX_RCA_ID_M11
  `undef AXI_MAX_RCA_ID_M11
`endif 

`ifdef AXI_LOG2_MAX_RCA_ID_P1_M11
  `undef AXI_LOG2_MAX_RCA_ID_P1_M11
`endif 

`ifdef AXI_MAX_WCA_ID_M11
  `undef AXI_MAX_WCA_ID_M11
`endif 

`ifdef AXI_LOG2_MAX_WCA_ID_P1_M11
  `undef AXI_LOG2_MAX_WCA_ID_P1_M11
`endif 

`ifdef AXI_MAX_URIDA_M11
  `undef AXI_MAX_URIDA_M11
`endif 

`ifdef AXI_LOG2_MAX_URIDA_M11
  `undef AXI_LOG2_MAX_URIDA_M11
`endif 

`ifdef AXI_MAX_UWIDA_M11
  `undef AXI_MAX_UWIDA_M11
`endif 

`ifdef AXI_LOG2_MAX_UWIDA_M11
  `undef AXI_LOG2_MAX_UWIDA_M11
`endif 

`ifdef AXI_RI_LIMIT_M11
  `undef AXI_RI_LIMIT_M11
`endif 

`ifdef AXI_MAX_RCA_ID_M12
  `undef AXI_MAX_RCA_ID_M12
`endif 

`ifdef AXI_LOG2_MAX_RCA_ID_P1_M12
  `undef AXI_LOG2_MAX_RCA_ID_P1_M12
`endif 

`ifdef AXI_MAX_WCA_ID_M12
  `undef AXI_MAX_WCA_ID_M12
`endif 

`ifdef AXI_LOG2_MAX_WCA_ID_P1_M12
  `undef AXI_LOG2_MAX_WCA_ID_P1_M12
`endif 

`ifdef AXI_MAX_URIDA_M12
  `undef AXI_MAX_URIDA_M12
`endif 

`ifdef AXI_LOG2_MAX_URIDA_M12
  `undef AXI_LOG2_MAX_URIDA_M12
`endif 

`ifdef AXI_MAX_UWIDA_M12
  `undef AXI_MAX_UWIDA_M12
`endif 

`ifdef AXI_LOG2_MAX_UWIDA_M12
  `undef AXI_LOG2_MAX_UWIDA_M12
`endif 

`ifdef AXI_RI_LIMIT_M12
  `undef AXI_RI_LIMIT_M12
`endif 

`ifdef AXI_MAX_RCA_ID_M13
  `undef AXI_MAX_RCA_ID_M13
`endif 

`ifdef AXI_LOG2_MAX_RCA_ID_P1_M13
  `undef AXI_LOG2_MAX_RCA_ID_P1_M13
`endif 

`ifdef AXI_MAX_WCA_ID_M13
  `undef AXI_MAX_WCA_ID_M13
`endif 

`ifdef AXI_LOG2_MAX_WCA_ID_P1_M13
  `undef AXI_LOG2_MAX_WCA_ID_P1_M13
`endif 

`ifdef AXI_MAX_URIDA_M13
  `undef AXI_MAX_URIDA_M13
`endif 

`ifdef AXI_LOG2_MAX_URIDA_M13
  `undef AXI_LOG2_MAX_URIDA_M13
`endif 

`ifdef AXI_MAX_UWIDA_M13
  `undef AXI_MAX_UWIDA_M13
`endif 

`ifdef AXI_LOG2_MAX_UWIDA_M13
  `undef AXI_LOG2_MAX_UWIDA_M13
`endif 

`ifdef AXI_RI_LIMIT_M13
  `undef AXI_RI_LIMIT_M13
`endif 

`ifdef AXI_MAX_RCA_ID_M14
  `undef AXI_MAX_RCA_ID_M14
`endif 

`ifdef AXI_LOG2_MAX_RCA_ID_P1_M14
  `undef AXI_LOG2_MAX_RCA_ID_P1_M14
`endif 

`ifdef AXI_MAX_WCA_ID_M14
  `undef AXI_MAX_WCA_ID_M14
`endif 

`ifdef AXI_LOG2_MAX_WCA_ID_P1_M14
  `undef AXI_LOG2_MAX_WCA_ID_P1_M14
`endif 

`ifdef AXI_MAX_URIDA_M14
  `undef AXI_MAX_URIDA_M14
`endif 

`ifdef AXI_LOG2_MAX_URIDA_M14
  `undef AXI_LOG2_MAX_URIDA_M14
`endif 

`ifdef AXI_MAX_UWIDA_M14
  `undef AXI_MAX_UWIDA_M14
`endif 

`ifdef AXI_LOG2_MAX_UWIDA_M14
  `undef AXI_LOG2_MAX_UWIDA_M14
`endif 

`ifdef AXI_RI_LIMIT_M14
  `undef AXI_RI_LIMIT_M14
`endif 

`ifdef AXI_MAX_RCA_ID_M15
  `undef AXI_MAX_RCA_ID_M15
`endif 

`ifdef AXI_LOG2_MAX_RCA_ID_P1_M15
  `undef AXI_LOG2_MAX_RCA_ID_P1_M15
`endif 

`ifdef AXI_MAX_WCA_ID_M15
  `undef AXI_MAX_WCA_ID_M15
`endif 

`ifdef AXI_LOG2_MAX_WCA_ID_P1_M15
  `undef AXI_LOG2_MAX_WCA_ID_P1_M15
`endif 

`ifdef AXI_MAX_URIDA_M15
  `undef AXI_MAX_URIDA_M15
`endif 

`ifdef AXI_LOG2_MAX_URIDA_M15
  `undef AXI_LOG2_MAX_URIDA_M15
`endif 

`ifdef AXI_MAX_UWIDA_M15
  `undef AXI_MAX_UWIDA_M15
`endif 

`ifdef AXI_LOG2_MAX_UWIDA_M15
  `undef AXI_LOG2_MAX_UWIDA_M15
`endif 

`ifdef AXI_RI_LIMIT_M15
  `undef AXI_RI_LIMIT_M15
`endif 

`ifdef AXI_MAX_RCA_ID_M16
  `undef AXI_MAX_RCA_ID_M16
`endif 

`ifdef AXI_LOG2_MAX_RCA_ID_P1_M16
  `undef AXI_LOG2_MAX_RCA_ID_P1_M16
`endif 

`ifdef AXI_MAX_WCA_ID_M16
  `undef AXI_MAX_WCA_ID_M16
`endif 

`ifdef AXI_LOG2_MAX_WCA_ID_P1_M16
  `undef AXI_LOG2_MAX_WCA_ID_P1_M16
`endif 

`ifdef AXI_MAX_URIDA_M16
  `undef AXI_MAX_URIDA_M16
`endif 

`ifdef AXI_LOG2_MAX_URIDA_M16
  `undef AXI_LOG2_MAX_URIDA_M16
`endif 

`ifdef AXI_MAX_UWIDA_M16
  `undef AXI_MAX_UWIDA_M16
`endif 

`ifdef AXI_LOG2_MAX_UWIDA_M16
  `undef AXI_LOG2_MAX_UWIDA_M16
`endif 

`ifdef AXI_RI_LIMIT_M16
  `undef AXI_RI_LIMIT_M16
`endif 

`ifdef AXI_MAX_FAWC_S0
  `undef AXI_MAX_FAWC_S0
`endif 

`ifdef AXI_LOG2_MAX_FAWC_S0
  `undef AXI_LOG2_MAX_FAWC_S0
`endif 

`ifdef AXI_LOG2_MAX_FAWC_P1_S0
  `undef AXI_LOG2_MAX_FAWC_P1_S0
`endif 

`ifdef AXI_MAX_FARC_S0
  `undef AXI_MAX_FARC_S0
`endif 

`ifdef AXI_LOG2_MAX_FARC_P1_S0
  `undef AXI_LOG2_MAX_FARC_P1_S0
`endif 

`ifdef AXI_WID_S0
  `undef AXI_WID_S0
`endif 

`ifdef AXI_MAX_FAC_EN
  `undef AXI_MAX_FAC_EN
`endif 

`ifdef AXI_WID_S1
  `undef AXI_WID_S1
`endif 

`ifdef AXI_LOG2_WID_S1
  `undef AXI_LOG2_WID_S1
`endif 

`ifdef AXI_LOG2_WID_P1_S1
  `undef AXI_LOG2_WID_P1_S1
`endif 

`ifdef AXI_MAX_FAWC_S1
  `undef AXI_MAX_FAWC_S1
`endif 

`ifdef AXI_LOG2_MAX_FAWC_S1
  `undef AXI_LOG2_MAX_FAWC_S1
`endif 

`ifdef AXI_LOG2_MAX_FAWC_P1_S1
  `undef AXI_LOG2_MAX_FAWC_P1_S1
`endif 

`ifdef AXI_MAX_FARC_S1
  `undef AXI_MAX_FARC_S1
`endif 

`ifdef AXI_LOG2_MAX_FARC_P1_S1
  `undef AXI_LOG2_MAX_FARC_P1_S1
`endif 

`ifdef AXI_WID_S2
  `undef AXI_WID_S2
`endif 

`ifdef AXI_LOG2_WID_S2
  `undef AXI_LOG2_WID_S2
`endif 

`ifdef AXI_LOG2_WID_P1_S2
  `undef AXI_LOG2_WID_P1_S2
`endif 

`ifdef AXI_MAX_FAWC_S2
  `undef AXI_MAX_FAWC_S2
`endif 

`ifdef AXI_LOG2_MAX_FAWC_S2
  `undef AXI_LOG2_MAX_FAWC_S2
`endif 

`ifdef AXI_LOG2_MAX_FAWC_P1_S2
  `undef AXI_LOG2_MAX_FAWC_P1_S2
`endif 

`ifdef AXI_MAX_FARC_S2
  `undef AXI_MAX_FARC_S2
`endif 

`ifdef AXI_LOG2_MAX_FARC_P1_S2
  `undef AXI_LOG2_MAX_FARC_P1_S2
`endif 

`ifdef AXI_WID_S3
  `undef AXI_WID_S3
`endif 

`ifdef AXI_LOG2_WID_S3
  `undef AXI_LOG2_WID_S3
`endif 

`ifdef AXI_LOG2_WID_P1_S3
  `undef AXI_LOG2_WID_P1_S3
`endif 

`ifdef AXI_MAX_FAWC_S3
  `undef AXI_MAX_FAWC_S3
`endif 

`ifdef AXI_LOG2_MAX_FAWC_S3
  `undef AXI_LOG2_MAX_FAWC_S3
`endif 

`ifdef AXI_LOG2_MAX_FAWC_P1_S3
  `undef AXI_LOG2_MAX_FAWC_P1_S3
`endif 

`ifdef AXI_MAX_FARC_S3
  `undef AXI_MAX_FARC_S3
`endif 

`ifdef AXI_LOG2_MAX_FARC_P1_S3
  `undef AXI_LOG2_MAX_FARC_P1_S3
`endif 

`ifdef AXI_WID_S4
  `undef AXI_WID_S4
`endif 

`ifdef AXI_LOG2_WID_S4
  `undef AXI_LOG2_WID_S4
`endif 

`ifdef AXI_LOG2_WID_P1_S4
  `undef AXI_LOG2_WID_P1_S4
`endif 

`ifdef AXI_MAX_FAWC_S4
  `undef AXI_MAX_FAWC_S4
`endif 

`ifdef AXI_LOG2_MAX_FAWC_S4
  `undef AXI_LOG2_MAX_FAWC_S4
`endif 

`ifdef AXI_LOG2_MAX_FAWC_P1_S4
  `undef AXI_LOG2_MAX_FAWC_P1_S4
`endif 

`ifdef AXI_MAX_FARC_S4
  `undef AXI_MAX_FARC_S4
`endif 

`ifdef AXI_LOG2_MAX_FARC_P1_S4
  `undef AXI_LOG2_MAX_FARC_P1_S4
`endif 

`ifdef AXI_WID_S5
  `undef AXI_WID_S5
`endif 

`ifdef AXI_LOG2_WID_S5
  `undef AXI_LOG2_WID_S5
`endif 

`ifdef AXI_LOG2_WID_P1_S5
  `undef AXI_LOG2_WID_P1_S5
`endif 

`ifdef AXI_MAX_FAWC_S5
  `undef AXI_MAX_FAWC_S5
`endif 

`ifdef AXI_LOG2_MAX_FAWC_S5
  `undef AXI_LOG2_MAX_FAWC_S5
`endif 

`ifdef AXI_LOG2_MAX_FAWC_P1_S5
  `undef AXI_LOG2_MAX_FAWC_P1_S5
`endif 

`ifdef AXI_MAX_FARC_S5
  `undef AXI_MAX_FARC_S5
`endif 

`ifdef AXI_LOG2_MAX_FARC_P1_S5
  `undef AXI_LOG2_MAX_FARC_P1_S5
`endif 

`ifdef AXI_WID_S6
  `undef AXI_WID_S6
`endif 

`ifdef AXI_LOG2_WID_S6
  `undef AXI_LOG2_WID_S6
`endif 

`ifdef AXI_LOG2_WID_P1_S6
  `undef AXI_LOG2_WID_P1_S6
`endif 

`ifdef AXI_MAX_FAWC_S6
  `undef AXI_MAX_FAWC_S6
`endif 

`ifdef AXI_LOG2_MAX_FAWC_S6
  `undef AXI_LOG2_MAX_FAWC_S6
`endif 

`ifdef AXI_LOG2_MAX_FAWC_P1_S6
  `undef AXI_LOG2_MAX_FAWC_P1_S6
`endif 

`ifdef AXI_MAX_FARC_S6
  `undef AXI_MAX_FARC_S6
`endif 

`ifdef AXI_LOG2_MAX_FARC_P1_S6
  `undef AXI_LOG2_MAX_FARC_P1_S6
`endif 

`ifdef AXI_WID_S7
  `undef AXI_WID_S7
`endif 

`ifdef AXI_LOG2_WID_S7
  `undef AXI_LOG2_WID_S7
`endif 

`ifdef AXI_LOG2_WID_P1_S7
  `undef AXI_LOG2_WID_P1_S7
`endif 

`ifdef AXI_MAX_FAWC_S7
  `undef AXI_MAX_FAWC_S7
`endif 

`ifdef AXI_LOG2_MAX_FAWC_S7
  `undef AXI_LOG2_MAX_FAWC_S7
`endif 

`ifdef AXI_LOG2_MAX_FAWC_P1_S7
  `undef AXI_LOG2_MAX_FAWC_P1_S7
`endif 

`ifdef AXI_MAX_FARC_S7
  `undef AXI_MAX_FARC_S7
`endif 

`ifdef AXI_LOG2_MAX_FARC_P1_S7
  `undef AXI_LOG2_MAX_FARC_P1_S7
`endif 

`ifdef AXI_WID_S8
  `undef AXI_WID_S8
`endif 

`ifdef AXI_LOG2_WID_S8
  `undef AXI_LOG2_WID_S8
`endif 

`ifdef AXI_LOG2_WID_P1_S8
  `undef AXI_LOG2_WID_P1_S8
`endif 

`ifdef AXI_MAX_FAWC_S8
  `undef AXI_MAX_FAWC_S8
`endif 

`ifdef AXI_LOG2_MAX_FAWC_S8
  `undef AXI_LOG2_MAX_FAWC_S8
`endif 

`ifdef AXI_LOG2_MAX_FAWC_P1_S8
  `undef AXI_LOG2_MAX_FAWC_P1_S8
`endif 

`ifdef AXI_MAX_FARC_S8
  `undef AXI_MAX_FARC_S8
`endif 

`ifdef AXI_LOG2_MAX_FARC_P1_S8
  `undef AXI_LOG2_MAX_FARC_P1_S8
`endif 

`ifdef AXI_WID_S9
  `undef AXI_WID_S9
`endif 

`ifdef AXI_LOG2_WID_S9
  `undef AXI_LOG2_WID_S9
`endif 

`ifdef AXI_LOG2_WID_P1_S9
  `undef AXI_LOG2_WID_P1_S9
`endif 

`ifdef AXI_MAX_FAWC_S9
  `undef AXI_MAX_FAWC_S9
`endif 

`ifdef AXI_LOG2_MAX_FAWC_S9
  `undef AXI_LOG2_MAX_FAWC_S9
`endif 

`ifdef AXI_LOG2_MAX_FAWC_P1_S9
  `undef AXI_LOG2_MAX_FAWC_P1_S9
`endif 

`ifdef AXI_MAX_FARC_S9
  `undef AXI_MAX_FARC_S9
`endif 

`ifdef AXI_LOG2_MAX_FARC_P1_S9
  `undef AXI_LOG2_MAX_FARC_P1_S9
`endif 

`ifdef AXI_WID_S10
  `undef AXI_WID_S10
`endif 

`ifdef AXI_LOG2_WID_S10
  `undef AXI_LOG2_WID_S10
`endif 

`ifdef AXI_LOG2_WID_P1_S10
  `undef AXI_LOG2_WID_P1_S10
`endif 

`ifdef AXI_MAX_FAWC_S10
  `undef AXI_MAX_FAWC_S10
`endif 

`ifdef AXI_LOG2_MAX_FAWC_S10
  `undef AXI_LOG2_MAX_FAWC_S10
`endif 

`ifdef AXI_LOG2_MAX_FAWC_P1_S10
  `undef AXI_LOG2_MAX_FAWC_P1_S10
`endif 

`ifdef AXI_MAX_FARC_S10
  `undef AXI_MAX_FARC_S10
`endif 

`ifdef AXI_LOG2_MAX_FARC_P1_S10
  `undef AXI_LOG2_MAX_FARC_P1_S10
`endif 

`ifdef AXI_WID_S11
  `undef AXI_WID_S11
`endif 

`ifdef AXI_LOG2_WID_S11
  `undef AXI_LOG2_WID_S11
`endif 

`ifdef AXI_LOG2_WID_P1_S11
  `undef AXI_LOG2_WID_P1_S11
`endif 

`ifdef AXI_MAX_FAWC_S11
  `undef AXI_MAX_FAWC_S11
`endif 

`ifdef AXI_LOG2_MAX_FAWC_S11
  `undef AXI_LOG2_MAX_FAWC_S11
`endif 

`ifdef AXI_LOG2_MAX_FAWC_P1_S11
  `undef AXI_LOG2_MAX_FAWC_P1_S11
`endif 

`ifdef AXI_MAX_FARC_S11
  `undef AXI_MAX_FARC_S11
`endif 

`ifdef AXI_LOG2_MAX_FARC_P1_S11
  `undef AXI_LOG2_MAX_FARC_P1_S11
`endif 

`ifdef AXI_WID_S12
  `undef AXI_WID_S12
`endif 

`ifdef AXI_LOG2_WID_S12
  `undef AXI_LOG2_WID_S12
`endif 

`ifdef AXI_LOG2_WID_P1_S12
  `undef AXI_LOG2_WID_P1_S12
`endif 

`ifdef AXI_MAX_FAWC_S12
  `undef AXI_MAX_FAWC_S12
`endif 

`ifdef AXI_LOG2_MAX_FAWC_S12
  `undef AXI_LOG2_MAX_FAWC_S12
`endif 

`ifdef AXI_LOG2_MAX_FAWC_P1_S12
  `undef AXI_LOG2_MAX_FAWC_P1_S12
`endif 

`ifdef AXI_MAX_FARC_S12
  `undef AXI_MAX_FARC_S12
`endif 

`ifdef AXI_LOG2_MAX_FARC_P1_S12
  `undef AXI_LOG2_MAX_FARC_P1_S12
`endif 

`ifdef AXI_WID_S13
  `undef AXI_WID_S13
`endif 

`ifdef AXI_LOG2_WID_S13
  `undef AXI_LOG2_WID_S13
`endif 

`ifdef AXI_LOG2_WID_P1_S13
  `undef AXI_LOG2_WID_P1_S13
`endif 

`ifdef AXI_MAX_FAWC_S13
  `undef AXI_MAX_FAWC_S13
`endif 

`ifdef AXI_LOG2_MAX_FAWC_S13
  `undef AXI_LOG2_MAX_FAWC_S13
`endif 

`ifdef AXI_LOG2_MAX_FAWC_P1_S13
  `undef AXI_LOG2_MAX_FAWC_P1_S13
`endif 

`ifdef AXI_MAX_FARC_S13
  `undef AXI_MAX_FARC_S13
`endif 

`ifdef AXI_LOG2_MAX_FARC_P1_S13
  `undef AXI_LOG2_MAX_FARC_P1_S13
`endif 

`ifdef AXI_WID_S14
  `undef AXI_WID_S14
`endif 

`ifdef AXI_LOG2_WID_S14
  `undef AXI_LOG2_WID_S14
`endif 

`ifdef AXI_LOG2_WID_P1_S14
  `undef AXI_LOG2_WID_P1_S14
`endif 

`ifdef AXI_MAX_FAWC_S14
  `undef AXI_MAX_FAWC_S14
`endif 

`ifdef AXI_LOG2_MAX_FAWC_S14
  `undef AXI_LOG2_MAX_FAWC_S14
`endif 

`ifdef AXI_LOG2_MAX_FAWC_P1_S14
  `undef AXI_LOG2_MAX_FAWC_P1_S14
`endif 

`ifdef AXI_MAX_FARC_S14
  `undef AXI_MAX_FARC_S14
`endif 

`ifdef AXI_LOG2_MAX_FARC_P1_S14
  `undef AXI_LOG2_MAX_FARC_P1_S14
`endif 

`ifdef AXI_WID_S15
  `undef AXI_WID_S15
`endif 

`ifdef AXI_LOG2_WID_S15
  `undef AXI_LOG2_WID_S15
`endif 

`ifdef AXI_LOG2_WID_P1_S15
  `undef AXI_LOG2_WID_P1_S15
`endif 

`ifdef AXI_MAX_FAWC_S15
  `undef AXI_MAX_FAWC_S15
`endif 

`ifdef AXI_LOG2_MAX_FAWC_S15
  `undef AXI_LOG2_MAX_FAWC_S15
`endif 

`ifdef AXI_LOG2_MAX_FAWC_P1_S15
  `undef AXI_LOG2_MAX_FAWC_P1_S15
`endif 

`ifdef AXI_MAX_FARC_S15
  `undef AXI_MAX_FARC_S15
`endif 

`ifdef AXI_LOG2_MAX_FARC_P1_S15
  `undef AXI_LOG2_MAX_FARC_P1_S15
`endif 

`ifdef AXI_WID_S16
  `undef AXI_WID_S16
`endif 

`ifdef AXI_LOG2_WID_S16
  `undef AXI_LOG2_WID_S16
`endif 

`ifdef AXI_LOG2_WID_P1_S16
  `undef AXI_LOG2_WID_P1_S16
`endif 

`ifdef AXI_MAX_FAWC_S16
  `undef AXI_MAX_FAWC_S16
`endif 

`ifdef AXI_LOG2_MAX_FAWC_S16
  `undef AXI_LOG2_MAX_FAWC_S16
`endif 

`ifdef AXI_LOG2_MAX_FAWC_P1_S16
  `undef AXI_LOG2_MAX_FAWC_P1_S16
`endif 

`ifdef AXI_MAX_FARC_S16
  `undef AXI_MAX_FARC_S16
`endif 

`ifdef AXI_LOG2_MAX_FARC_P1_S16
  `undef AXI_LOG2_MAX_FARC_P1_S16
`endif 

`ifdef AXI_S0_SHARED_FARC
  `undef AXI_S0_SHARED_FARC
`endif 

`ifdef AXI_LOG2_S0_SHARED_FARC_P1
  `undef AXI_LOG2_S0_SHARED_FARC_P1
`endif 

`ifdef AXI_S0_SHARED_AR_HAS_DDCTD
  `undef AXI_S0_SHARED_AR_HAS_DDCTD
`endif 

`ifdef AXI_S0_SHARED_FAWC
  `undef AXI_S0_SHARED_FAWC
`endif 

`ifdef AXI_LOG2_S0_SHARED_FAWC_P1
  `undef AXI_LOG2_S0_SHARED_FAWC_P1
`endif 

`ifdef AXI_S0_SHARED_AW_HAS_DDCTD
  `undef AXI_S0_SHARED_AW_HAS_DDCTD
`endif 

`ifdef AXI_S0_SHARED_W_HAS_DDCTD
  `undef AXI_S0_SHARED_W_HAS_DDCTD
`endif 

`ifdef AXI_S1_SHARED_FARC
  `undef AXI_S1_SHARED_FARC
`endif 

`ifdef AXI_LOG2_S1_SHARED_FARC_P1
  `undef AXI_LOG2_S1_SHARED_FARC_P1
`endif 

`ifdef AXI_S1_SHARED_AR_HAS_DDCTD
  `undef AXI_S1_SHARED_AR_HAS_DDCTD
`endif 

`ifdef AXI_S1_SHARED_FAWC
  `undef AXI_S1_SHARED_FAWC
`endif 

`ifdef AXI_LOG2_S1_SHARED_FAWC_P1
  `undef AXI_LOG2_S1_SHARED_FAWC_P1
`endif 

`ifdef AXI_S1_SHARED_AW_HAS_DDCTD
  `undef AXI_S1_SHARED_AW_HAS_DDCTD
`endif 

`ifdef AXI_S1_SHARED_W_HAS_DDCTD
  `undef AXI_S1_SHARED_W_HAS_DDCTD
`endif 

`ifdef AXI_S2_SHARED_FARC
  `undef AXI_S2_SHARED_FARC
`endif 

`ifdef AXI_LOG2_S2_SHARED_FARC_P1
  `undef AXI_LOG2_S2_SHARED_FARC_P1
`endif 

`ifdef AXI_S2_SHARED_AR_HAS_DDCTD
  `undef AXI_S2_SHARED_AR_HAS_DDCTD
`endif 

`ifdef AXI_S2_SHARED_FAWC
  `undef AXI_S2_SHARED_FAWC
`endif 

`ifdef AXI_LOG2_S2_SHARED_FAWC_P1
  `undef AXI_LOG2_S2_SHARED_FAWC_P1
`endif 

`ifdef AXI_S2_SHARED_AW_HAS_DDCTD
  `undef AXI_S2_SHARED_AW_HAS_DDCTD
`endif 

`ifdef AXI_S2_SHARED_W_HAS_DDCTD
  `undef AXI_S2_SHARED_W_HAS_DDCTD
`endif 

`ifdef AXI_S3_SHARED_FARC
  `undef AXI_S3_SHARED_FARC
`endif 

`ifdef AXI_LOG2_S3_SHARED_FARC_P1
  `undef AXI_LOG2_S3_SHARED_FARC_P1
`endif 

`ifdef AXI_S3_SHARED_AR_HAS_DDCTD
  `undef AXI_S3_SHARED_AR_HAS_DDCTD
`endif 

`ifdef AXI_S3_SHARED_FAWC
  `undef AXI_S3_SHARED_FAWC
`endif 

`ifdef AXI_LOG2_S3_SHARED_FAWC_P1
  `undef AXI_LOG2_S3_SHARED_FAWC_P1
`endif 

`ifdef AXI_S3_SHARED_AW_HAS_DDCTD
  `undef AXI_S3_SHARED_AW_HAS_DDCTD
`endif 

`ifdef AXI_S3_SHARED_W_HAS_DDCTD
  `undef AXI_S3_SHARED_W_HAS_DDCTD
`endif 

`ifdef AXI_S4_SHARED_FARC
  `undef AXI_S4_SHARED_FARC
`endif 

`ifdef AXI_LOG2_S4_SHARED_FARC_P1
  `undef AXI_LOG2_S4_SHARED_FARC_P1
`endif 

`ifdef AXI_S4_SHARED_AR_HAS_DDCTD
  `undef AXI_S4_SHARED_AR_HAS_DDCTD
`endif 

`ifdef AXI_S4_SHARED_FAWC
  `undef AXI_S4_SHARED_FAWC
`endif 

`ifdef AXI_LOG2_S4_SHARED_FAWC_P1
  `undef AXI_LOG2_S4_SHARED_FAWC_P1
`endif 

`ifdef AXI_S4_SHARED_AW_HAS_DDCTD
  `undef AXI_S4_SHARED_AW_HAS_DDCTD
`endif 

`ifdef AXI_S4_SHARED_W_HAS_DDCTD
  `undef AXI_S4_SHARED_W_HAS_DDCTD
`endif 

`ifdef AXI_S5_SHARED_FARC
  `undef AXI_S5_SHARED_FARC
`endif 

`ifdef AXI_LOG2_S5_SHARED_FARC_P1
  `undef AXI_LOG2_S5_SHARED_FARC_P1
`endif 

`ifdef AXI_S5_SHARED_AR_HAS_DDCTD
  `undef AXI_S5_SHARED_AR_HAS_DDCTD
`endif 

`ifdef AXI_S5_SHARED_FAWC
  `undef AXI_S5_SHARED_FAWC
`endif 

`ifdef AXI_LOG2_S5_SHARED_FAWC_P1
  `undef AXI_LOG2_S5_SHARED_FAWC_P1
`endif 

`ifdef AXI_S5_SHARED_AW_HAS_DDCTD
  `undef AXI_S5_SHARED_AW_HAS_DDCTD
`endif 

`ifdef AXI_S5_SHARED_W_HAS_DDCTD
  `undef AXI_S5_SHARED_W_HAS_DDCTD
`endif 

`ifdef AXI_S6_SHARED_FARC
  `undef AXI_S6_SHARED_FARC
`endif 

`ifdef AXI_LOG2_S6_SHARED_FARC_P1
  `undef AXI_LOG2_S6_SHARED_FARC_P1
`endif 

`ifdef AXI_S6_SHARED_AR_HAS_DDCTD
  `undef AXI_S6_SHARED_AR_HAS_DDCTD
`endif 

`ifdef AXI_S6_SHARED_FAWC
  `undef AXI_S6_SHARED_FAWC
`endif 

`ifdef AXI_LOG2_S6_SHARED_FAWC_P1
  `undef AXI_LOG2_S6_SHARED_FAWC_P1
`endif 

`ifdef AXI_S6_SHARED_AW_HAS_DDCTD
  `undef AXI_S6_SHARED_AW_HAS_DDCTD
`endif 

`ifdef AXI_S6_SHARED_W_HAS_DDCTD
  `undef AXI_S6_SHARED_W_HAS_DDCTD
`endif 

`ifdef AXI_S7_SHARED_FARC
  `undef AXI_S7_SHARED_FARC
`endif 

`ifdef AXI_LOG2_S7_SHARED_FARC_P1
  `undef AXI_LOG2_S7_SHARED_FARC_P1
`endif 

`ifdef AXI_S7_SHARED_AR_HAS_DDCTD
  `undef AXI_S7_SHARED_AR_HAS_DDCTD
`endif 

`ifdef AXI_S7_SHARED_FAWC
  `undef AXI_S7_SHARED_FAWC
`endif 

`ifdef AXI_LOG2_S7_SHARED_FAWC_P1
  `undef AXI_LOG2_S7_SHARED_FAWC_P1
`endif 

`ifdef AXI_S7_SHARED_AW_HAS_DDCTD
  `undef AXI_S7_SHARED_AW_HAS_DDCTD
`endif 

`ifdef AXI_S7_SHARED_W_HAS_DDCTD
  `undef AXI_S7_SHARED_W_HAS_DDCTD
`endif 

`ifdef AXI_S8_SHARED_FARC
  `undef AXI_S8_SHARED_FARC
`endif 

`ifdef AXI_LOG2_S8_SHARED_FARC_P1
  `undef AXI_LOG2_S8_SHARED_FARC_P1
`endif 

`ifdef AXI_S8_SHARED_AR_HAS_DDCTD
  `undef AXI_S8_SHARED_AR_HAS_DDCTD
`endif 

`ifdef AXI_S8_SHARED_FAWC
  `undef AXI_S8_SHARED_FAWC
`endif 

`ifdef AXI_LOG2_S8_SHARED_FAWC_P1
  `undef AXI_LOG2_S8_SHARED_FAWC_P1
`endif 

`ifdef AXI_S8_SHARED_AW_HAS_DDCTD
  `undef AXI_S8_SHARED_AW_HAS_DDCTD
`endif 

`ifdef AXI_S8_SHARED_W_HAS_DDCTD
  `undef AXI_S8_SHARED_W_HAS_DDCTD
`endif 

`ifdef AXI_S9_SHARED_FARC
  `undef AXI_S9_SHARED_FARC
`endif 

`ifdef AXI_LOG2_S9_SHARED_FARC_P1
  `undef AXI_LOG2_S9_SHARED_FARC_P1
`endif 

`ifdef AXI_S9_SHARED_AR_HAS_DDCTD
  `undef AXI_S9_SHARED_AR_HAS_DDCTD
`endif 

`ifdef AXI_S9_SHARED_FAWC
  `undef AXI_S9_SHARED_FAWC
`endif 

`ifdef AXI_LOG2_S9_SHARED_FAWC_P1
  `undef AXI_LOG2_S9_SHARED_FAWC_P1
`endif 

`ifdef AXI_S9_SHARED_AW_HAS_DDCTD
  `undef AXI_S9_SHARED_AW_HAS_DDCTD
`endif 

`ifdef AXI_S9_SHARED_W_HAS_DDCTD
  `undef AXI_S9_SHARED_W_HAS_DDCTD
`endif 

`ifdef AXI_S10_SHARED_FARC
  `undef AXI_S10_SHARED_FARC
`endif 

`ifdef AXI_LOG2_S10_SHARED_FARC_P1
  `undef AXI_LOG2_S10_SHARED_FARC_P1
`endif 

`ifdef AXI_S10_SHARED_AR_HAS_DDCTD
  `undef AXI_S10_SHARED_AR_HAS_DDCTD
`endif 

`ifdef AXI_S10_SHARED_FAWC
  `undef AXI_S10_SHARED_FAWC
`endif 

`ifdef AXI_LOG2_S10_SHARED_FAWC_P1
  `undef AXI_LOG2_S10_SHARED_FAWC_P1
`endif 

`ifdef AXI_S10_SHARED_AW_HAS_DDCTD
  `undef AXI_S10_SHARED_AW_HAS_DDCTD
`endif 

`ifdef AXI_S10_SHARED_W_HAS_DDCTD
  `undef AXI_S10_SHARED_W_HAS_DDCTD
`endif 

`ifdef AXI_S11_SHARED_FARC
  `undef AXI_S11_SHARED_FARC
`endif 

`ifdef AXI_LOG2_S11_SHARED_FARC_P1
  `undef AXI_LOG2_S11_SHARED_FARC_P1
`endif 

`ifdef AXI_S11_SHARED_AR_HAS_DDCTD
  `undef AXI_S11_SHARED_AR_HAS_DDCTD
`endif 

`ifdef AXI_S11_SHARED_FAWC
  `undef AXI_S11_SHARED_FAWC
`endif 

`ifdef AXI_LOG2_S11_SHARED_FAWC_P1
  `undef AXI_LOG2_S11_SHARED_FAWC_P1
`endif 

`ifdef AXI_S11_SHARED_AW_HAS_DDCTD
  `undef AXI_S11_SHARED_AW_HAS_DDCTD
`endif 

`ifdef AXI_S11_SHARED_W_HAS_DDCTD
  `undef AXI_S11_SHARED_W_HAS_DDCTD
`endif 

`ifdef AXI_S12_SHARED_FARC
  `undef AXI_S12_SHARED_FARC
`endif 

`ifdef AXI_LOG2_S12_SHARED_FARC_P1
  `undef AXI_LOG2_S12_SHARED_FARC_P1
`endif 

`ifdef AXI_S12_SHARED_AR_HAS_DDCTD
  `undef AXI_S12_SHARED_AR_HAS_DDCTD
`endif 

`ifdef AXI_S12_SHARED_FAWC
  `undef AXI_S12_SHARED_FAWC
`endif 

`ifdef AXI_LOG2_S12_SHARED_FAWC_P1
  `undef AXI_LOG2_S12_SHARED_FAWC_P1
`endif 

`ifdef AXI_S12_SHARED_AW_HAS_DDCTD
  `undef AXI_S12_SHARED_AW_HAS_DDCTD
`endif 

`ifdef AXI_S12_SHARED_W_HAS_DDCTD
  `undef AXI_S12_SHARED_W_HAS_DDCTD
`endif 

`ifdef AXI_S13_SHARED_FARC
  `undef AXI_S13_SHARED_FARC
`endif 

`ifdef AXI_LOG2_S13_SHARED_FARC_P1
  `undef AXI_LOG2_S13_SHARED_FARC_P1
`endif 

`ifdef AXI_S13_SHARED_AR_HAS_DDCTD
  `undef AXI_S13_SHARED_AR_HAS_DDCTD
`endif 

`ifdef AXI_S13_SHARED_FAWC
  `undef AXI_S13_SHARED_FAWC
`endif 

`ifdef AXI_LOG2_S13_SHARED_FAWC_P1
  `undef AXI_LOG2_S13_SHARED_FAWC_P1
`endif 

`ifdef AXI_S13_SHARED_AW_HAS_DDCTD
  `undef AXI_S13_SHARED_AW_HAS_DDCTD
`endif 

`ifdef AXI_S13_SHARED_W_HAS_DDCTD
  `undef AXI_S13_SHARED_W_HAS_DDCTD
`endif 

`ifdef AXI_S14_SHARED_FARC
  `undef AXI_S14_SHARED_FARC
`endif 

`ifdef AXI_LOG2_S14_SHARED_FARC_P1
  `undef AXI_LOG2_S14_SHARED_FARC_P1
`endif 

`ifdef AXI_S14_SHARED_AR_HAS_DDCTD
  `undef AXI_S14_SHARED_AR_HAS_DDCTD
`endif 

`ifdef AXI_S14_SHARED_FAWC
  `undef AXI_S14_SHARED_FAWC
`endif 

`ifdef AXI_LOG2_S14_SHARED_FAWC_P1
  `undef AXI_LOG2_S14_SHARED_FAWC_P1
`endif 

`ifdef AXI_S14_SHARED_AW_HAS_DDCTD
  `undef AXI_S14_SHARED_AW_HAS_DDCTD
`endif 

`ifdef AXI_S14_SHARED_W_HAS_DDCTD
  `undef AXI_S14_SHARED_W_HAS_DDCTD
`endif 

`ifdef AXI_S15_SHARED_FARC
  `undef AXI_S15_SHARED_FARC
`endif 

`ifdef AXI_LOG2_S15_SHARED_FARC_P1
  `undef AXI_LOG2_S15_SHARED_FARC_P1
`endif 

`ifdef AXI_S15_SHARED_AR_HAS_DDCTD
  `undef AXI_S15_SHARED_AR_HAS_DDCTD
`endif 

`ifdef AXI_S15_SHARED_FAWC
  `undef AXI_S15_SHARED_FAWC
`endif 

`ifdef AXI_LOG2_S15_SHARED_FAWC_P1
  `undef AXI_LOG2_S15_SHARED_FAWC_P1
`endif 

`ifdef AXI_S15_SHARED_AW_HAS_DDCTD
  `undef AXI_S15_SHARED_AW_HAS_DDCTD
`endif 

`ifdef AXI_S15_SHARED_W_HAS_DDCTD
  `undef AXI_S15_SHARED_W_HAS_DDCTD
`endif 

`ifdef AXI_S16_SHARED_FARC
  `undef AXI_S16_SHARED_FARC
`endif 

`ifdef AXI_LOG2_S16_SHARED_FARC_P1
  `undef AXI_LOG2_S16_SHARED_FARC_P1
`endif 

`ifdef AXI_S16_SHARED_AR_HAS_DDCTD
  `undef AXI_S16_SHARED_AR_HAS_DDCTD
`endif 

`ifdef AXI_S16_SHARED_FAWC
  `undef AXI_S16_SHARED_FAWC
`endif 

`ifdef AXI_LOG2_S16_SHARED_FAWC_P1
  `undef AXI_LOG2_S16_SHARED_FAWC_P1
`endif 

`ifdef AXI_S16_SHARED_AW_HAS_DDCTD
  `undef AXI_S16_SHARED_AW_HAS_DDCTD
`endif 

`ifdef AXI_S16_SHARED_W_HAS_DDCTD
  `undef AXI_S16_SHARED_W_HAS_DDCTD
`endif 

`ifdef AXI_M0_SHARED_R_HAS_DDCTD
  `undef AXI_M0_SHARED_R_HAS_DDCTD
`endif 

`ifdef AXI_M0_SHARED_B_HAS_DDCTD
  `undef AXI_M0_SHARED_B_HAS_DDCTD
`endif 

`ifdef AXI_M1_SHARED_R_HAS_DDCTD
  `undef AXI_M1_SHARED_R_HAS_DDCTD
`endif 

`ifdef AXI_M1_SHARED_B_HAS_DDCTD
  `undef AXI_M1_SHARED_B_HAS_DDCTD
`endif 

`ifdef AXI_M2_SHARED_R_HAS_DDCTD
  `undef AXI_M2_SHARED_R_HAS_DDCTD
`endif 

`ifdef AXI_M2_SHARED_B_HAS_DDCTD
  `undef AXI_M2_SHARED_B_HAS_DDCTD
`endif 

`ifdef AXI_M3_SHARED_R_HAS_DDCTD
  `undef AXI_M3_SHARED_R_HAS_DDCTD
`endif 

`ifdef AXI_M3_SHARED_B_HAS_DDCTD
  `undef AXI_M3_SHARED_B_HAS_DDCTD
`endif 

`ifdef AXI_M4_SHARED_R_HAS_DDCTD
  `undef AXI_M4_SHARED_R_HAS_DDCTD
`endif 

`ifdef AXI_M4_SHARED_B_HAS_DDCTD
  `undef AXI_M4_SHARED_B_HAS_DDCTD
`endif 

`ifdef AXI_M5_SHARED_R_HAS_DDCTD
  `undef AXI_M5_SHARED_R_HAS_DDCTD
`endif 

`ifdef AXI_M5_SHARED_B_HAS_DDCTD
  `undef AXI_M5_SHARED_B_HAS_DDCTD
`endif 

`ifdef AXI_M6_SHARED_R_HAS_DDCTD
  `undef AXI_M6_SHARED_R_HAS_DDCTD
`endif 

`ifdef AXI_M6_SHARED_B_HAS_DDCTD
  `undef AXI_M6_SHARED_B_HAS_DDCTD
`endif 

`ifdef AXI_M7_SHARED_R_HAS_DDCTD
  `undef AXI_M7_SHARED_R_HAS_DDCTD
`endif 

`ifdef AXI_M7_SHARED_B_HAS_DDCTD
  `undef AXI_M7_SHARED_B_HAS_DDCTD
`endif 

`ifdef AXI_M8_SHARED_R_HAS_DDCTD
  `undef AXI_M8_SHARED_R_HAS_DDCTD
`endif 

`ifdef AXI_M8_SHARED_B_HAS_DDCTD
  `undef AXI_M8_SHARED_B_HAS_DDCTD
`endif 

`ifdef AXI_M9_SHARED_R_HAS_DDCTD
  `undef AXI_M9_SHARED_R_HAS_DDCTD
`endif 

`ifdef AXI_M9_SHARED_B_HAS_DDCTD
  `undef AXI_M9_SHARED_B_HAS_DDCTD
`endif 

`ifdef AXI_M10_SHARED_R_HAS_DDCTD
  `undef AXI_M10_SHARED_R_HAS_DDCTD
`endif 

`ifdef AXI_M10_SHARED_B_HAS_DDCTD
  `undef AXI_M10_SHARED_B_HAS_DDCTD
`endif 

`ifdef AXI_M11_SHARED_R_HAS_DDCTD
  `undef AXI_M11_SHARED_R_HAS_DDCTD
`endif 

`ifdef AXI_M11_SHARED_B_HAS_DDCTD
  `undef AXI_M11_SHARED_B_HAS_DDCTD
`endif 

`ifdef AXI_M12_SHARED_R_HAS_DDCTD
  `undef AXI_M12_SHARED_R_HAS_DDCTD
`endif 

`ifdef AXI_M12_SHARED_B_HAS_DDCTD
  `undef AXI_M12_SHARED_B_HAS_DDCTD
`endif 

`ifdef AXI_M13_SHARED_R_HAS_DDCTD
  `undef AXI_M13_SHARED_R_HAS_DDCTD
`endif 

`ifdef AXI_M13_SHARED_B_HAS_DDCTD
  `undef AXI_M13_SHARED_B_HAS_DDCTD
`endif 

`ifdef AXI_M14_SHARED_R_HAS_DDCTD
  `undef AXI_M14_SHARED_R_HAS_DDCTD
`endif 

`ifdef AXI_M14_SHARED_B_HAS_DDCTD
  `undef AXI_M14_SHARED_B_HAS_DDCTD
`endif 

`ifdef AXI_M15_SHARED_R_HAS_DDCTD
  `undef AXI_M15_SHARED_R_HAS_DDCTD
`endif 

`ifdef AXI_M15_SHARED_B_HAS_DDCTD
  `undef AXI_M15_SHARED_B_HAS_DDCTD
`endif 

`ifdef AXI_PRIORITY_M1
  `undef AXI_PRIORITY_M1
`endif 

`ifdef AXI_PRIORITY_M2
  `undef AXI_PRIORITY_M2
`endif 

`ifdef AXI_PRIORITY_M3
  `undef AXI_PRIORITY_M3
`endif 

`ifdef AXI_PRIORITY_M4
  `undef AXI_PRIORITY_M4
`endif 

`ifdef AXI_PRIORITY_M5
  `undef AXI_PRIORITY_M5
`endif 

`ifdef AXI_PRIORITY_M6
  `undef AXI_PRIORITY_M6
`endif 

`ifdef AXI_PRIORITY_M7
  `undef AXI_PRIORITY_M7
`endif 

`ifdef AXI_PRIORITY_M8
  `undef AXI_PRIORITY_M8
`endif 

`ifdef AXI_PRIORITY_M9
  `undef AXI_PRIORITY_M9
`endif 

`ifdef AXI_PRIORITY_M10
  `undef AXI_PRIORITY_M10
`endif 

`ifdef AXI_PRIORITY_M11
  `undef AXI_PRIORITY_M11
`endif 

`ifdef AXI_PRIORITY_M12
  `undef AXI_PRIORITY_M12
`endif 

`ifdef AXI_PRIORITY_M13
  `undef AXI_PRIORITY_M13
`endif 

`ifdef AXI_PRIORITY_M14
  `undef AXI_PRIORITY_M14
`endif 

`ifdef AXI_PRIORITY_M15
  `undef AXI_PRIORITY_M15
`endif 

`ifdef AXI_PRIORITY_M16
  `undef AXI_PRIORITY_M16
`endif 

`ifdef AXI_PRIORITY_S1
  `undef AXI_PRIORITY_S1
`endif 

`ifdef AXI_PRIORITY_S2
  `undef AXI_PRIORITY_S2
`endif 

`ifdef AXI_PRIORITY_S3
  `undef AXI_PRIORITY_S3
`endif 

`ifdef AXI_PRIORITY_S4
  `undef AXI_PRIORITY_S4
`endif 

`ifdef AXI_PRIORITY_S5
  `undef AXI_PRIORITY_S5
`endif 

`ifdef AXI_PRIORITY_S6
  `undef AXI_PRIORITY_S6
`endif 

`ifdef AXI_PRIORITY_S7
  `undef AXI_PRIORITY_S7
`endif 

`ifdef AXI_PRIORITY_S8
  `undef AXI_PRIORITY_S8
`endif 

`ifdef AXI_PRIORITY_S9
  `undef AXI_PRIORITY_S9
`endif 

`ifdef AXI_PRIORITY_S10
  `undef AXI_PRIORITY_S10
`endif 

`ifdef AXI_PRIORITY_S11
  `undef AXI_PRIORITY_S11
`endif 

`ifdef AXI_PRIORITY_S12
  `undef AXI_PRIORITY_S12
`endif 

`ifdef AXI_PRIORITY_S13
  `undef AXI_PRIORITY_S13
`endif 

`ifdef AXI_PRIORITY_S14
  `undef AXI_PRIORITY_S14
`endif 

`ifdef AXI_PRIORITY_S15
  `undef AXI_PRIORITY_S15
`endif 

`ifdef AXI_PRIORITY_S16
  `undef AXI_PRIORITY_S16
`endif 

`ifdef AXI_PRIORITY_S0
  `undef AXI_PRIORITY_S0
`endif 

`ifdef AXI_HAS_EXT_PRIORITY
  `undef AXI_HAS_EXT_PRIORITY
`endif 

`ifdef AXI_SHARED_LAYER_MASTER_PRIORITY_EN_VAL
  `undef AXI_SHARED_LAYER_MASTER_PRIORITY_EN_VAL
`endif 

`ifdef AXI_SHARED_LAYER_MASTER_PRIORITY_EN
  `undef AXI_SHARED_LAYER_MASTER_PRIORITY_EN
`endif 

`ifdef AXI_SHARED_LAYER_MASTER_PRIORITY
  `undef AXI_SHARED_LAYER_MASTER_PRIORITY
`endif 

`ifdef AXI_SHARED_LAYER_SLAVE_PRIORITY_EN_VAL
  `undef AXI_SHARED_LAYER_SLAVE_PRIORITY_EN_VAL
`endif 

`ifdef AXI_SHARED_LAYER_SLAVE_PRIORITY_EN
  `undef AXI_SHARED_LAYER_SLAVE_PRIORITY_EN
`endif 

`ifdef AXI_SHARED_LAYER_SLAVE_PRIORITY
  `undef AXI_SHARED_LAYER_SLAVE_PRIORITY
`endif 

`ifdef AXI_AR_ARB_TYPE_S0
  `undef AXI_AR_ARB_TYPE_S0
`endif 

`ifdef AXI_AW_ARB_TYPE_S0
  `undef AXI_AW_ARB_TYPE_S0
`endif 

`ifdef AXI_AR_ARB_TYPE_S1
  `undef AXI_AR_ARB_TYPE_S1
`endif 

`ifdef AXI_AW_ARB_TYPE_S1
  `undef AXI_AW_ARB_TYPE_S1
`endif 

`ifdef AXI_AR_ARB_TYPE_S2
  `undef AXI_AR_ARB_TYPE_S2
`endif 

`ifdef AXI_AW_ARB_TYPE_S2
  `undef AXI_AW_ARB_TYPE_S2
`endif 

`ifdef AXI_AR_ARB_TYPE_S3
  `undef AXI_AR_ARB_TYPE_S3
`endif 

`ifdef AXI_AW_ARB_TYPE_S3
  `undef AXI_AW_ARB_TYPE_S3
`endif 

`ifdef AXI_AR_ARB_TYPE_S4
  `undef AXI_AR_ARB_TYPE_S4
`endif 

`ifdef AXI_AW_ARB_TYPE_S4
  `undef AXI_AW_ARB_TYPE_S4
`endif 

`ifdef AXI_AR_ARB_TYPE_S5
  `undef AXI_AR_ARB_TYPE_S5
`endif 

`ifdef AXI_AW_ARB_TYPE_S5
  `undef AXI_AW_ARB_TYPE_S5
`endif 

`ifdef AXI_AR_ARB_TYPE_S6
  `undef AXI_AR_ARB_TYPE_S6
`endif 

`ifdef AXI_AW_ARB_TYPE_S6
  `undef AXI_AW_ARB_TYPE_S6
`endif 

`ifdef AXI_AR_ARB_TYPE_S7
  `undef AXI_AR_ARB_TYPE_S7
`endif 

`ifdef AXI_AW_ARB_TYPE_S7
  `undef AXI_AW_ARB_TYPE_S7
`endif 

`ifdef AXI_AR_ARB_TYPE_S8
  `undef AXI_AR_ARB_TYPE_S8
`endif 

`ifdef AXI_AW_ARB_TYPE_S8
  `undef AXI_AW_ARB_TYPE_S8
`endif 

`ifdef AXI_AR_ARB_TYPE_S9
  `undef AXI_AR_ARB_TYPE_S9
`endif 

`ifdef AXI_AW_ARB_TYPE_S9
  `undef AXI_AW_ARB_TYPE_S9
`endif 

`ifdef AXI_AR_ARB_TYPE_S10
  `undef AXI_AR_ARB_TYPE_S10
`endif 

`ifdef AXI_AW_ARB_TYPE_S10
  `undef AXI_AW_ARB_TYPE_S10
`endif 

`ifdef AXI_AR_ARB_TYPE_S11
  `undef AXI_AR_ARB_TYPE_S11
`endif 

`ifdef AXI_AW_ARB_TYPE_S11
  `undef AXI_AW_ARB_TYPE_S11
`endif 

`ifdef AXI_AR_ARB_TYPE_S12
  `undef AXI_AR_ARB_TYPE_S12
`endif 

`ifdef AXI_AW_ARB_TYPE_S12
  `undef AXI_AW_ARB_TYPE_S12
`endif 

`ifdef AXI_AR_ARB_TYPE_S13
  `undef AXI_AR_ARB_TYPE_S13
`endif 

`ifdef AXI_AW_ARB_TYPE_S13
  `undef AXI_AW_ARB_TYPE_S13
`endif 

`ifdef AXI_AR_ARB_TYPE_S14
  `undef AXI_AR_ARB_TYPE_S14
`endif 

`ifdef AXI_AW_ARB_TYPE_S14
  `undef AXI_AW_ARB_TYPE_S14
`endif 

`ifdef AXI_AR_ARB_TYPE_S15
  `undef AXI_AR_ARB_TYPE_S15
`endif 

`ifdef AXI_AW_ARB_TYPE_S15
  `undef AXI_AW_ARB_TYPE_S15
`endif 

`ifdef AXI_AR_ARB_TYPE_S16
  `undef AXI_AR_ARB_TYPE_S16
`endif 

`ifdef AXI_AW_ARB_TYPE_S16
  `undef AXI_AW_ARB_TYPE_S16
`endif 

`ifdef AXI_W_ARB_TYPE_S0
  `undef AXI_W_ARB_TYPE_S0
`endif 

`ifdef AXI_W_ARB_TYPE_S1
  `undef AXI_W_ARB_TYPE_S1
`endif 

`ifdef AXI_W_ARB_TYPE_S2
  `undef AXI_W_ARB_TYPE_S2
`endif 

`ifdef AXI_W_ARB_TYPE_S3
  `undef AXI_W_ARB_TYPE_S3
`endif 

`ifdef AXI_W_ARB_TYPE_S4
  `undef AXI_W_ARB_TYPE_S4
`endif 

`ifdef AXI_W_ARB_TYPE_S5
  `undef AXI_W_ARB_TYPE_S5
`endif 

`ifdef AXI_W_ARB_TYPE_S6
  `undef AXI_W_ARB_TYPE_S6
`endif 

`ifdef AXI_W_ARB_TYPE_S7
  `undef AXI_W_ARB_TYPE_S7
`endif 

`ifdef AXI_W_ARB_TYPE_S8
  `undef AXI_W_ARB_TYPE_S8
`endif 

`ifdef AXI_W_ARB_TYPE_S9
  `undef AXI_W_ARB_TYPE_S9
`endif 

`ifdef AXI_W_ARB_TYPE_S10
  `undef AXI_W_ARB_TYPE_S10
`endif 

`ifdef AXI_W_ARB_TYPE_S11
  `undef AXI_W_ARB_TYPE_S11
`endif 

`ifdef AXI_W_ARB_TYPE_S12
  `undef AXI_W_ARB_TYPE_S12
`endif 

`ifdef AXI_W_ARB_TYPE_S13
  `undef AXI_W_ARB_TYPE_S13
`endif 

`ifdef AXI_W_ARB_TYPE_S14
  `undef AXI_W_ARB_TYPE_S14
`endif 

`ifdef AXI_W_ARB_TYPE_S15
  `undef AXI_W_ARB_TYPE_S15
`endif 

`ifdef AXI_W_ARB_TYPE_S16
  `undef AXI_W_ARB_TYPE_S16
`endif 

`ifdef AXI_R_ARB_TYPE_M1
  `undef AXI_R_ARB_TYPE_M1
`endif 

`ifdef AXI_B_ARB_TYPE_M1
  `undef AXI_B_ARB_TYPE_M1
`endif 

`ifdef AXI_R_ARB_TYPE_M2
  `undef AXI_R_ARB_TYPE_M2
`endif 

`ifdef AXI_B_ARB_TYPE_M2
  `undef AXI_B_ARB_TYPE_M2
`endif 

`ifdef AXI_R_ARB_TYPE_M3
  `undef AXI_R_ARB_TYPE_M3
`endif 

`ifdef AXI_B_ARB_TYPE_M3
  `undef AXI_B_ARB_TYPE_M3
`endif 

`ifdef AXI_R_ARB_TYPE_M4
  `undef AXI_R_ARB_TYPE_M4
`endif 

`ifdef AXI_B_ARB_TYPE_M4
  `undef AXI_B_ARB_TYPE_M4
`endif 

`ifdef AXI_R_ARB_TYPE_M5
  `undef AXI_R_ARB_TYPE_M5
`endif 

`ifdef AXI_B_ARB_TYPE_M5
  `undef AXI_B_ARB_TYPE_M5
`endif 

`ifdef AXI_R_ARB_TYPE_M6
  `undef AXI_R_ARB_TYPE_M6
`endif 

`ifdef AXI_B_ARB_TYPE_M6
  `undef AXI_B_ARB_TYPE_M6
`endif 

`ifdef AXI_R_ARB_TYPE_M7
  `undef AXI_R_ARB_TYPE_M7
`endif 

`ifdef AXI_B_ARB_TYPE_M7
  `undef AXI_B_ARB_TYPE_M7
`endif 

`ifdef AXI_R_ARB_TYPE_M8
  `undef AXI_R_ARB_TYPE_M8
`endif 

`ifdef AXI_B_ARB_TYPE_M8
  `undef AXI_B_ARB_TYPE_M8
`endif 

`ifdef AXI_R_ARB_TYPE_M9
  `undef AXI_R_ARB_TYPE_M9
`endif 

`ifdef AXI_B_ARB_TYPE_M9
  `undef AXI_B_ARB_TYPE_M9
`endif 

`ifdef AXI_R_ARB_TYPE_M10
  `undef AXI_R_ARB_TYPE_M10
`endif 

`ifdef AXI_B_ARB_TYPE_M10
  `undef AXI_B_ARB_TYPE_M10
`endif 

`ifdef AXI_R_ARB_TYPE_M11
  `undef AXI_R_ARB_TYPE_M11
`endif 

`ifdef AXI_B_ARB_TYPE_M11
  `undef AXI_B_ARB_TYPE_M11
`endif 

`ifdef AXI_R_ARB_TYPE_M12
  `undef AXI_R_ARB_TYPE_M12
`endif 

`ifdef AXI_B_ARB_TYPE_M12
  `undef AXI_B_ARB_TYPE_M12
`endif 

`ifdef AXI_R_ARB_TYPE_M13
  `undef AXI_R_ARB_TYPE_M13
`endif 

`ifdef AXI_B_ARB_TYPE_M13
  `undef AXI_B_ARB_TYPE_M13
`endif 

`ifdef AXI_R_ARB_TYPE_M14
  `undef AXI_R_ARB_TYPE_M14
`endif 

`ifdef AXI_B_ARB_TYPE_M14
  `undef AXI_B_ARB_TYPE_M14
`endif 

`ifdef AXI_R_ARB_TYPE_M15
  `undef AXI_R_ARB_TYPE_M15
`endif 

`ifdef AXI_B_ARB_TYPE_M15
  `undef AXI_B_ARB_TYPE_M15
`endif 

`ifdef AXI_R_ARB_TYPE_M16
  `undef AXI_R_ARB_TYPE_M16
`endif 

`ifdef AXI_B_ARB_TYPE_M16
  `undef AXI_B_ARB_TYPE_M16
`endif 

`ifdef AXI_AR_SHARED_ARB_TYPE
  `undef AXI_AR_SHARED_ARB_TYPE
`endif 

`ifdef AXI_AW_SHARED_ARB_TYPE
  `undef AXI_AW_SHARED_ARB_TYPE
`endif 

`ifdef AXI_W_SHARED_ARB_TYPE
  `undef AXI_W_SHARED_ARB_TYPE
`endif 

`ifdef AXI_R_SHARED_ARB_TYPE
  `undef AXI_R_SHARED_ARB_TYPE
`endif 

`ifdef AXI_B_SHARED_ARB_TYPE
  `undef AXI_B_SHARED_ARB_TYPE
`endif 

`ifdef AXI_USER_ARB_REMOVAL
  `undef AXI_USER_ARB_REMOVAL
`endif 

`ifdef AXI_NUM_RN_S1
  `undef AXI_NUM_RN_S1
`endif 

`ifdef AXI_NUM_RN_S2
  `undef AXI_NUM_RN_S2
`endif 

`ifdef AXI_NUM_RN_S3
  `undef AXI_NUM_RN_S3
`endif 

`ifdef AXI_NUM_RN_S4
  `undef AXI_NUM_RN_S4
`endif 

`ifdef AXI_NUM_RN_S5
  `undef AXI_NUM_RN_S5
`endif 

`ifdef AXI_NUM_RN_S6
  `undef AXI_NUM_RN_S6
`endif 

`ifdef AXI_NUM_RN_S7
  `undef AXI_NUM_RN_S7
`endif 

`ifdef AXI_NUM_RN_S8
  `undef AXI_NUM_RN_S8
`endif 

`ifdef AXI_NUM_RN_S9
  `undef AXI_NUM_RN_S9
`endif 

`ifdef AXI_NUM_RN_S10
  `undef AXI_NUM_RN_S10
`endif 

`ifdef AXI_NUM_RN_S11
  `undef AXI_NUM_RN_S11
`endif 

`ifdef AXI_NUM_RN_S12
  `undef AXI_NUM_RN_S12
`endif 

`ifdef AXI_NUM_RN_S13
  `undef AXI_NUM_RN_S13
`endif 

`ifdef AXI_NUM_RN_S14
  `undef AXI_NUM_RN_S14
`endif 

`ifdef AXI_NUM_RN_S15
  `undef AXI_NUM_RN_S15
`endif 

`ifdef AXI_NUM_RN_S16
  `undef AXI_NUM_RN_S16
`endif 

`ifdef AXI_R1_NSA_S1
  `undef AXI_R1_NSA_S1
`endif 

`ifdef AXI_R1_NEA_S1
  `undef AXI_R1_NEA_S1
`endif 

`ifdef AXI_R1_NSA_S2
  `undef AXI_R1_NSA_S2
`endif 

`ifdef AXI_R1_NEA_S2
  `undef AXI_R1_NEA_S2
`endif 

`ifdef AXI_R1_NSA_S3
  `undef AXI_R1_NSA_S3
`endif 

`ifdef AXI_R1_NEA_S3
  `undef AXI_R1_NEA_S3
`endif 

`ifdef AXI_R1_NSA_S4
  `undef AXI_R1_NSA_S4
`endif 

`ifdef AXI_R1_NEA_S4
  `undef AXI_R1_NEA_S4
`endif 

`ifdef AXI_R1_NSA_S5
  `undef AXI_R1_NSA_S5
`endif 

`ifdef AXI_R1_NEA_S5
  `undef AXI_R1_NEA_S5
`endif 

`ifdef AXI_R1_NSA_S6
  `undef AXI_R1_NSA_S6
`endif 

`ifdef AXI_R1_NEA_S6
  `undef AXI_R1_NEA_S6
`endif 

`ifdef AXI_R1_NSA_S7
  `undef AXI_R1_NSA_S7
`endif 

`ifdef AXI_R1_NEA_S7
  `undef AXI_R1_NEA_S7
`endif 

`ifdef AXI_R1_NSA_S8
  `undef AXI_R1_NSA_S8
`endif 

`ifdef AXI_R1_NEA_S8
  `undef AXI_R1_NEA_S8
`endif 

`ifdef AXI_R1_NSA_S9
  `undef AXI_R1_NSA_S9
`endif 

`ifdef AXI_R1_NEA_S9
  `undef AXI_R1_NEA_S9
`endif 

`ifdef AXI_R1_NSA_S10
  `undef AXI_R1_NSA_S10
`endif 

`ifdef AXI_R1_NEA_S10
  `undef AXI_R1_NEA_S10
`endif 

`ifdef AXI_R1_NSA_S11
  `undef AXI_R1_NSA_S11
`endif 

`ifdef AXI_R1_NEA_S11
  `undef AXI_R1_NEA_S11
`endif 

`ifdef AXI_R1_NSA_S12
  `undef AXI_R1_NSA_S12
`endif 

`ifdef AXI_R1_NEA_S12
  `undef AXI_R1_NEA_S12
`endif 

`ifdef AXI_R1_NSA_S13
  `undef AXI_R1_NSA_S13
`endif 

`ifdef AXI_R1_NEA_S13
  `undef AXI_R1_NEA_S13
`endif 

`ifdef AXI_R1_NSA_S14
  `undef AXI_R1_NSA_S14
`endif 

`ifdef AXI_R1_NEA_S14
  `undef AXI_R1_NEA_S14
`endif 

`ifdef AXI_R1_NSA_S15
  `undef AXI_R1_NSA_S15
`endif 

`ifdef AXI_R1_NEA_S15
  `undef AXI_R1_NEA_S15
`endif 

`ifdef AXI_R1_NSA_S16
  `undef AXI_R1_NSA_S16
`endif 

`ifdef AXI_R1_NEA_S16
  `undef AXI_R1_NEA_S16
`endif 

`ifdef AXI_R2_NSA_S1
  `undef AXI_R2_NSA_S1
`endif 

`ifdef AXI_R2_NEA_S1
  `undef AXI_R2_NEA_S1
`endif 

`ifdef AXI_R2_NSA_S2
  `undef AXI_R2_NSA_S2
`endif 

`ifdef AXI_R2_NEA_S2
  `undef AXI_R2_NEA_S2
`endif 

`ifdef AXI_R2_NSA_S3
  `undef AXI_R2_NSA_S3
`endif 

`ifdef AXI_R2_NEA_S3
  `undef AXI_R2_NEA_S3
`endif 

`ifdef AXI_R2_NSA_S4
  `undef AXI_R2_NSA_S4
`endif 

`ifdef AXI_R2_NEA_S4
  `undef AXI_R2_NEA_S4
`endif 

`ifdef AXI_R2_NSA_S5
  `undef AXI_R2_NSA_S5
`endif 

`ifdef AXI_R2_NEA_S5
  `undef AXI_R2_NEA_S5
`endif 

`ifdef AXI_R2_NSA_S6
  `undef AXI_R2_NSA_S6
`endif 

`ifdef AXI_R2_NEA_S6
  `undef AXI_R2_NEA_S6
`endif 

`ifdef AXI_R2_NSA_S7
  `undef AXI_R2_NSA_S7
`endif 

`ifdef AXI_R2_NEA_S7
  `undef AXI_R2_NEA_S7
`endif 

`ifdef AXI_R2_NSA_S8
  `undef AXI_R2_NSA_S8
`endif 

`ifdef AXI_R2_NEA_S8
  `undef AXI_R2_NEA_S8
`endif 

`ifdef AXI_R2_NSA_S9
  `undef AXI_R2_NSA_S9
`endif 

`ifdef AXI_R2_NEA_S9
  `undef AXI_R2_NEA_S9
`endif 

`ifdef AXI_R2_NSA_S10
  `undef AXI_R2_NSA_S10
`endif 

`ifdef AXI_R2_NEA_S10
  `undef AXI_R2_NEA_S10
`endif 

`ifdef AXI_R2_NSA_S11
  `undef AXI_R2_NSA_S11
`endif 

`ifdef AXI_R2_NEA_S11
  `undef AXI_R2_NEA_S11
`endif 

`ifdef AXI_R2_NSA_S12
  `undef AXI_R2_NSA_S12
`endif 

`ifdef AXI_R2_NEA_S12
  `undef AXI_R2_NEA_S12
`endif 

`ifdef AXI_R2_NSA_S13
  `undef AXI_R2_NSA_S13
`endif 

`ifdef AXI_R2_NEA_S13
  `undef AXI_R2_NEA_S13
`endif 

`ifdef AXI_R2_NSA_S14
  `undef AXI_R2_NSA_S14
`endif 

`ifdef AXI_R2_NEA_S14
  `undef AXI_R2_NEA_S14
`endif 

`ifdef AXI_R2_NSA_S15
  `undef AXI_R2_NSA_S15
`endif 

`ifdef AXI_R2_NEA_S15
  `undef AXI_R2_NEA_S15
`endif 

`ifdef AXI_R2_NSA_S16
  `undef AXI_R2_NSA_S16
`endif 

`ifdef AXI_R2_NEA_S16
  `undef AXI_R2_NEA_S16
`endif 

`ifdef AXI_R3_NSA_S1
  `undef AXI_R3_NSA_S1
`endif 

`ifdef AXI_R3_NEA_S1
  `undef AXI_R3_NEA_S1
`endif 

`ifdef AXI_R3_NSA_S2
  `undef AXI_R3_NSA_S2
`endif 

`ifdef AXI_R3_NEA_S2
  `undef AXI_R3_NEA_S2
`endif 

`ifdef AXI_R3_NSA_S3
  `undef AXI_R3_NSA_S3
`endif 

`ifdef AXI_R3_NEA_S3
  `undef AXI_R3_NEA_S3
`endif 

`ifdef AXI_R3_NSA_S4
  `undef AXI_R3_NSA_S4
`endif 

`ifdef AXI_R3_NEA_S4
  `undef AXI_R3_NEA_S4
`endif 

`ifdef AXI_R3_NSA_S5
  `undef AXI_R3_NSA_S5
`endif 

`ifdef AXI_R3_NEA_S5
  `undef AXI_R3_NEA_S5
`endif 

`ifdef AXI_R3_NSA_S6
  `undef AXI_R3_NSA_S6
`endif 

`ifdef AXI_R3_NEA_S6
  `undef AXI_R3_NEA_S6
`endif 

`ifdef AXI_R3_NSA_S7
  `undef AXI_R3_NSA_S7
`endif 

`ifdef AXI_R3_NEA_S7
  `undef AXI_R3_NEA_S7
`endif 

`ifdef AXI_R3_NSA_S8
  `undef AXI_R3_NSA_S8
`endif 

`ifdef AXI_R3_NEA_S8
  `undef AXI_R3_NEA_S8
`endif 

`ifdef AXI_R3_NSA_S9
  `undef AXI_R3_NSA_S9
`endif 

`ifdef AXI_R3_NEA_S9
  `undef AXI_R3_NEA_S9
`endif 

`ifdef AXI_R3_NSA_S10
  `undef AXI_R3_NSA_S10
`endif 

`ifdef AXI_R3_NEA_S10
  `undef AXI_R3_NEA_S10
`endif 

`ifdef AXI_R3_NSA_S11
  `undef AXI_R3_NSA_S11
`endif 

`ifdef AXI_R3_NEA_S11
  `undef AXI_R3_NEA_S11
`endif 

`ifdef AXI_R3_NSA_S12
  `undef AXI_R3_NSA_S12
`endif 

`ifdef AXI_R3_NEA_S12
  `undef AXI_R3_NEA_S12
`endif 

`ifdef AXI_R3_NSA_S13
  `undef AXI_R3_NSA_S13
`endif 

`ifdef AXI_R3_NEA_S13
  `undef AXI_R3_NEA_S13
`endif 

`ifdef AXI_R3_NSA_S14
  `undef AXI_R3_NSA_S14
`endif 

`ifdef AXI_R3_NEA_S14
  `undef AXI_R3_NEA_S14
`endif 

`ifdef AXI_R3_NSA_S15
  `undef AXI_R3_NSA_S15
`endif 

`ifdef AXI_R3_NEA_S15
  `undef AXI_R3_NEA_S15
`endif 

`ifdef AXI_R3_NSA_S16
  `undef AXI_R3_NSA_S16
`endif 

`ifdef AXI_R3_NEA_S16
  `undef AXI_R3_NEA_S16
`endif 

`ifdef AXI_R4_NSA_S1
  `undef AXI_R4_NSA_S1
`endif 

`ifdef AXI_R4_NEA_S1
  `undef AXI_R4_NEA_S1
`endif 

`ifdef AXI_R4_NSA_S2
  `undef AXI_R4_NSA_S2
`endif 

`ifdef AXI_R4_NEA_S2
  `undef AXI_R4_NEA_S2
`endif 

`ifdef AXI_R4_NSA_S3
  `undef AXI_R4_NSA_S3
`endif 

`ifdef AXI_R4_NEA_S3
  `undef AXI_R4_NEA_S3
`endif 

`ifdef AXI_R4_NSA_S4
  `undef AXI_R4_NSA_S4
`endif 

`ifdef AXI_R4_NEA_S4
  `undef AXI_R4_NEA_S4
`endif 

`ifdef AXI_R4_NSA_S5
  `undef AXI_R4_NSA_S5
`endif 

`ifdef AXI_R4_NEA_S5
  `undef AXI_R4_NEA_S5
`endif 

`ifdef AXI_R4_NSA_S6
  `undef AXI_R4_NSA_S6
`endif 

`ifdef AXI_R4_NEA_S6
  `undef AXI_R4_NEA_S6
`endif 

`ifdef AXI_R4_NSA_S7
  `undef AXI_R4_NSA_S7
`endif 

`ifdef AXI_R4_NEA_S7
  `undef AXI_R4_NEA_S7
`endif 

`ifdef AXI_R4_NSA_S8
  `undef AXI_R4_NSA_S8
`endif 

`ifdef AXI_R4_NEA_S8
  `undef AXI_R4_NEA_S8
`endif 

`ifdef AXI_R4_NSA_S9
  `undef AXI_R4_NSA_S9
`endif 

`ifdef AXI_R4_NEA_S9
  `undef AXI_R4_NEA_S9
`endif 

`ifdef AXI_R4_NSA_S10
  `undef AXI_R4_NSA_S10
`endif 

`ifdef AXI_R4_NEA_S10
  `undef AXI_R4_NEA_S10
`endif 

`ifdef AXI_R4_NSA_S11
  `undef AXI_R4_NSA_S11
`endif 

`ifdef AXI_R4_NEA_S11
  `undef AXI_R4_NEA_S11
`endif 

`ifdef AXI_R4_NSA_S12
  `undef AXI_R4_NSA_S12
`endif 

`ifdef AXI_R4_NEA_S12
  `undef AXI_R4_NEA_S12
`endif 

`ifdef AXI_R4_NSA_S13
  `undef AXI_R4_NSA_S13
`endif 

`ifdef AXI_R4_NEA_S13
  `undef AXI_R4_NEA_S13
`endif 

`ifdef AXI_R4_NSA_S14
  `undef AXI_R4_NSA_S14
`endif 

`ifdef AXI_R4_NEA_S14
  `undef AXI_R4_NEA_S14
`endif 

`ifdef AXI_R4_NSA_S15
  `undef AXI_R4_NSA_S15
`endif 

`ifdef AXI_R4_NEA_S15
  `undef AXI_R4_NEA_S15
`endif 

`ifdef AXI_R4_NSA_S16
  `undef AXI_R4_NSA_S16
`endif 

`ifdef AXI_R4_NEA_S16
  `undef AXI_R4_NEA_S16
`endif 

`ifdef AXI_R5_NSA_S1
  `undef AXI_R5_NSA_S1
`endif 

`ifdef AXI_R5_NEA_S1
  `undef AXI_R5_NEA_S1
`endif 

`ifdef AXI_R5_NSA_S2
  `undef AXI_R5_NSA_S2
`endif 

`ifdef AXI_R5_NEA_S2
  `undef AXI_R5_NEA_S2
`endif 

`ifdef AXI_R5_NSA_S3
  `undef AXI_R5_NSA_S3
`endif 

`ifdef AXI_R5_NEA_S3
  `undef AXI_R5_NEA_S3
`endif 

`ifdef AXI_R5_NSA_S4
  `undef AXI_R5_NSA_S4
`endif 

`ifdef AXI_R5_NEA_S4
  `undef AXI_R5_NEA_S4
`endif 

`ifdef AXI_R5_NSA_S5
  `undef AXI_R5_NSA_S5
`endif 

`ifdef AXI_R5_NEA_S5
  `undef AXI_R5_NEA_S5
`endif 

`ifdef AXI_R5_NSA_S6
  `undef AXI_R5_NSA_S6
`endif 

`ifdef AXI_R5_NEA_S6
  `undef AXI_R5_NEA_S6
`endif 

`ifdef AXI_R5_NSA_S7
  `undef AXI_R5_NSA_S7
`endif 

`ifdef AXI_R5_NEA_S7
  `undef AXI_R5_NEA_S7
`endif 

`ifdef AXI_R5_NSA_S8
  `undef AXI_R5_NSA_S8
`endif 

`ifdef AXI_R5_NEA_S8
  `undef AXI_R5_NEA_S8
`endif 

`ifdef AXI_R5_NSA_S9
  `undef AXI_R5_NSA_S9
`endif 

`ifdef AXI_R5_NEA_S9
  `undef AXI_R5_NEA_S9
`endif 

`ifdef AXI_R5_NSA_S10
  `undef AXI_R5_NSA_S10
`endif 

`ifdef AXI_R5_NEA_S10
  `undef AXI_R5_NEA_S10
`endif 

`ifdef AXI_R5_NSA_S11
  `undef AXI_R5_NSA_S11
`endif 

`ifdef AXI_R5_NEA_S11
  `undef AXI_R5_NEA_S11
`endif 

`ifdef AXI_R5_NSA_S12
  `undef AXI_R5_NSA_S12
`endif 

`ifdef AXI_R5_NEA_S12
  `undef AXI_R5_NEA_S12
`endif 

`ifdef AXI_R5_NSA_S13
  `undef AXI_R5_NSA_S13
`endif 

`ifdef AXI_R5_NEA_S13
  `undef AXI_R5_NEA_S13
`endif 

`ifdef AXI_R5_NSA_S14
  `undef AXI_R5_NSA_S14
`endif 

`ifdef AXI_R5_NEA_S14
  `undef AXI_R5_NEA_S14
`endif 

`ifdef AXI_R5_NSA_S15
  `undef AXI_R5_NSA_S15
`endif 

`ifdef AXI_R5_NEA_S15
  `undef AXI_R5_NEA_S15
`endif 

`ifdef AXI_R5_NSA_S16
  `undef AXI_R5_NSA_S16
`endif 

`ifdef AXI_R5_NEA_S16
  `undef AXI_R5_NEA_S16
`endif 

`ifdef AXI_R6_NSA_S1
  `undef AXI_R6_NSA_S1
`endif 

`ifdef AXI_R6_NEA_S1
  `undef AXI_R6_NEA_S1
`endif 

`ifdef AXI_R6_NSA_S2
  `undef AXI_R6_NSA_S2
`endif 

`ifdef AXI_R6_NEA_S2
  `undef AXI_R6_NEA_S2
`endif 

`ifdef AXI_R6_NSA_S3
  `undef AXI_R6_NSA_S3
`endif 

`ifdef AXI_R6_NEA_S3
  `undef AXI_R6_NEA_S3
`endif 

`ifdef AXI_R6_NSA_S4
  `undef AXI_R6_NSA_S4
`endif 

`ifdef AXI_R6_NEA_S4
  `undef AXI_R6_NEA_S4
`endif 

`ifdef AXI_R6_NSA_S5
  `undef AXI_R6_NSA_S5
`endif 

`ifdef AXI_R6_NEA_S5
  `undef AXI_R6_NEA_S5
`endif 

`ifdef AXI_R6_NSA_S6
  `undef AXI_R6_NSA_S6
`endif 

`ifdef AXI_R6_NEA_S6
  `undef AXI_R6_NEA_S6
`endif 

`ifdef AXI_R6_NSA_S7
  `undef AXI_R6_NSA_S7
`endif 

`ifdef AXI_R6_NEA_S7
  `undef AXI_R6_NEA_S7
`endif 

`ifdef AXI_R6_NSA_S8
  `undef AXI_R6_NSA_S8
`endif 

`ifdef AXI_R6_NEA_S8
  `undef AXI_R6_NEA_S8
`endif 

`ifdef AXI_R6_NSA_S9
  `undef AXI_R6_NSA_S9
`endif 

`ifdef AXI_R6_NEA_S9
  `undef AXI_R6_NEA_S9
`endif 

`ifdef AXI_R6_NSA_S10
  `undef AXI_R6_NSA_S10
`endif 

`ifdef AXI_R6_NEA_S10
  `undef AXI_R6_NEA_S10
`endif 

`ifdef AXI_R6_NSA_S11
  `undef AXI_R6_NSA_S11
`endif 

`ifdef AXI_R6_NEA_S11
  `undef AXI_R6_NEA_S11
`endif 

`ifdef AXI_R6_NSA_S12
  `undef AXI_R6_NSA_S12
`endif 

`ifdef AXI_R6_NEA_S12
  `undef AXI_R6_NEA_S12
`endif 

`ifdef AXI_R6_NSA_S13
  `undef AXI_R6_NSA_S13
`endif 

`ifdef AXI_R6_NEA_S13
  `undef AXI_R6_NEA_S13
`endif 

`ifdef AXI_R6_NSA_S14
  `undef AXI_R6_NSA_S14
`endif 

`ifdef AXI_R6_NEA_S14
  `undef AXI_R6_NEA_S14
`endif 

`ifdef AXI_R6_NSA_S15
  `undef AXI_R6_NSA_S15
`endif 

`ifdef AXI_R6_NEA_S15
  `undef AXI_R6_NEA_S15
`endif 

`ifdef AXI_R6_NSA_S16
  `undef AXI_R6_NSA_S16
`endif 

`ifdef AXI_R6_NEA_S16
  `undef AXI_R6_NEA_S16
`endif 

`ifdef AXI_R7_NSA_S1
  `undef AXI_R7_NSA_S1
`endif 

`ifdef AXI_R7_NEA_S1
  `undef AXI_R7_NEA_S1
`endif 

`ifdef AXI_R7_NSA_S2
  `undef AXI_R7_NSA_S2
`endif 

`ifdef AXI_R7_NEA_S2
  `undef AXI_R7_NEA_S2
`endif 

`ifdef AXI_R7_NSA_S3
  `undef AXI_R7_NSA_S3
`endif 

`ifdef AXI_R7_NEA_S3
  `undef AXI_R7_NEA_S3
`endif 

`ifdef AXI_R7_NSA_S4
  `undef AXI_R7_NSA_S4
`endif 

`ifdef AXI_R7_NEA_S4
  `undef AXI_R7_NEA_S4
`endif 

`ifdef AXI_R7_NSA_S5
  `undef AXI_R7_NSA_S5
`endif 

`ifdef AXI_R7_NEA_S5
  `undef AXI_R7_NEA_S5
`endif 

`ifdef AXI_R7_NSA_S6
  `undef AXI_R7_NSA_S6
`endif 

`ifdef AXI_R7_NEA_S6
  `undef AXI_R7_NEA_S6
`endif 

`ifdef AXI_R7_NSA_S7
  `undef AXI_R7_NSA_S7
`endif 

`ifdef AXI_R7_NEA_S7
  `undef AXI_R7_NEA_S7
`endif 

`ifdef AXI_R7_NSA_S8
  `undef AXI_R7_NSA_S8
`endif 

`ifdef AXI_R7_NEA_S8
  `undef AXI_R7_NEA_S8
`endif 

`ifdef AXI_R7_NSA_S9
  `undef AXI_R7_NSA_S9
`endif 

`ifdef AXI_R7_NEA_S9
  `undef AXI_R7_NEA_S9
`endif 

`ifdef AXI_R7_NSA_S10
  `undef AXI_R7_NSA_S10
`endif 

`ifdef AXI_R7_NEA_S10
  `undef AXI_R7_NEA_S10
`endif 

`ifdef AXI_R7_NSA_S11
  `undef AXI_R7_NSA_S11
`endif 

`ifdef AXI_R7_NEA_S11
  `undef AXI_R7_NEA_S11
`endif 

`ifdef AXI_R7_NSA_S12
  `undef AXI_R7_NSA_S12
`endif 

`ifdef AXI_R7_NEA_S12
  `undef AXI_R7_NEA_S12
`endif 

`ifdef AXI_R7_NSA_S13
  `undef AXI_R7_NSA_S13
`endif 

`ifdef AXI_R7_NEA_S13
  `undef AXI_R7_NEA_S13
`endif 

`ifdef AXI_R7_NSA_S14
  `undef AXI_R7_NSA_S14
`endif 

`ifdef AXI_R7_NEA_S14
  `undef AXI_R7_NEA_S14
`endif 

`ifdef AXI_R7_NSA_S15
  `undef AXI_R7_NSA_S15
`endif 

`ifdef AXI_R7_NEA_S15
  `undef AXI_R7_NEA_S15
`endif 

`ifdef AXI_R7_NSA_S16
  `undef AXI_R7_NSA_S16
`endif 

`ifdef AXI_R7_NEA_S16
  `undef AXI_R7_NEA_S16
`endif 

`ifdef AXI_R8_NSA_S1
  `undef AXI_R8_NSA_S1
`endif 

`ifdef AXI_R8_NEA_S1
  `undef AXI_R8_NEA_S1
`endif 

`ifdef AXI_R8_NSA_S2
  `undef AXI_R8_NSA_S2
`endif 

`ifdef AXI_R8_NEA_S2
  `undef AXI_R8_NEA_S2
`endif 

`ifdef AXI_R8_NSA_S3
  `undef AXI_R8_NSA_S3
`endif 

`ifdef AXI_R8_NEA_S3
  `undef AXI_R8_NEA_S3
`endif 

`ifdef AXI_R8_NSA_S4
  `undef AXI_R8_NSA_S4
`endif 

`ifdef AXI_R8_NEA_S4
  `undef AXI_R8_NEA_S4
`endif 

`ifdef AXI_R8_NSA_S5
  `undef AXI_R8_NSA_S5
`endif 

`ifdef AXI_R8_NEA_S5
  `undef AXI_R8_NEA_S5
`endif 

`ifdef AXI_R8_NSA_S6
  `undef AXI_R8_NSA_S6
`endif 

`ifdef AXI_R8_NEA_S6
  `undef AXI_R8_NEA_S6
`endif 

`ifdef AXI_R8_NSA_S7
  `undef AXI_R8_NSA_S7
`endif 

`ifdef AXI_R8_NEA_S7
  `undef AXI_R8_NEA_S7
`endif 

`ifdef AXI_R8_NSA_S8
  `undef AXI_R8_NSA_S8
`endif 

`ifdef AXI_R8_NEA_S8
  `undef AXI_R8_NEA_S8
`endif 

`ifdef AXI_R8_NSA_S9
  `undef AXI_R8_NSA_S9
`endif 

`ifdef AXI_R8_NEA_S9
  `undef AXI_R8_NEA_S9
`endif 

`ifdef AXI_R8_NSA_S10
  `undef AXI_R8_NSA_S10
`endif 

`ifdef AXI_R8_NEA_S10
  `undef AXI_R8_NEA_S10
`endif 

`ifdef AXI_R8_NSA_S11
  `undef AXI_R8_NSA_S11
`endif 

`ifdef AXI_R8_NEA_S11
  `undef AXI_R8_NEA_S11
`endif 

`ifdef AXI_R8_NSA_S12
  `undef AXI_R8_NSA_S12
`endif 

`ifdef AXI_R8_NEA_S12
  `undef AXI_R8_NEA_S12
`endif 

`ifdef AXI_R8_NSA_S13
  `undef AXI_R8_NSA_S13
`endif 

`ifdef AXI_R8_NEA_S13
  `undef AXI_R8_NEA_S13
`endif 

`ifdef AXI_R8_NSA_S14
  `undef AXI_R8_NSA_S14
`endif 

`ifdef AXI_R8_NEA_S14
  `undef AXI_R8_NEA_S14
`endif 

`ifdef AXI_R8_NSA_S15
  `undef AXI_R8_NSA_S15
`endif 

`ifdef AXI_R8_NEA_S15
  `undef AXI_R8_NEA_S15
`endif 

`ifdef AXI_R8_NSA_S16
  `undef AXI_R8_NSA_S16
`endif 

`ifdef AXI_R8_NEA_S16
  `undef AXI_R8_NEA_S16
`endif 

`ifdef AXI_NUM_RB_S1
  `undef AXI_NUM_RB_S1
`endif 

`ifdef AXI_NUM_RB_S2
  `undef AXI_NUM_RB_S2
`endif 

`ifdef AXI_NUM_RB_S3
  `undef AXI_NUM_RB_S3
`endif 

`ifdef AXI_NUM_RB_S4
  `undef AXI_NUM_RB_S4
`endif 

`ifdef AXI_NUM_RB_S5
  `undef AXI_NUM_RB_S5
`endif 

`ifdef AXI_NUM_RB_S6
  `undef AXI_NUM_RB_S6
`endif 

`ifdef AXI_NUM_RB_S7
  `undef AXI_NUM_RB_S7
`endif 

`ifdef AXI_NUM_RB_S8
  `undef AXI_NUM_RB_S8
`endif 

`ifdef AXI_NUM_RB_S9
  `undef AXI_NUM_RB_S9
`endif 

`ifdef AXI_NUM_RB_S10
  `undef AXI_NUM_RB_S10
`endif 

`ifdef AXI_NUM_RB_S11
  `undef AXI_NUM_RB_S11
`endif 

`ifdef AXI_NUM_RB_S12
  `undef AXI_NUM_RB_S12
`endif 

`ifdef AXI_NUM_RB_S13
  `undef AXI_NUM_RB_S13
`endif 

`ifdef AXI_NUM_RB_S14
  `undef AXI_NUM_RB_S14
`endif 

`ifdef AXI_NUM_RB_S15
  `undef AXI_NUM_RB_S15
`endif 

`ifdef AXI_NUM_RB_S16
  `undef AXI_NUM_RB_S16
`endif 

`ifdef AXI_R1_BSA_S1
  `undef AXI_R1_BSA_S1
`endif 

`ifdef AXI_R1_BEA_S1
  `undef AXI_R1_BEA_S1
`endif 

`ifdef AXI_R1_BSA_S2
  `undef AXI_R1_BSA_S2
`endif 

`ifdef AXI_R1_BEA_S2
  `undef AXI_R1_BEA_S2
`endif 

`ifdef AXI_R1_BSA_S3
  `undef AXI_R1_BSA_S3
`endif 

`ifdef AXI_R1_BEA_S3
  `undef AXI_R1_BEA_S3
`endif 

`ifdef AXI_R1_BSA_S4
  `undef AXI_R1_BSA_S4
`endif 

`ifdef AXI_R1_BEA_S4
  `undef AXI_R1_BEA_S4
`endif 

`ifdef AXI_R1_BSA_S5
  `undef AXI_R1_BSA_S5
`endif 

`ifdef AXI_R1_BEA_S5
  `undef AXI_R1_BEA_S5
`endif 

`ifdef AXI_R1_BSA_S6
  `undef AXI_R1_BSA_S6
`endif 

`ifdef AXI_R1_BEA_S6
  `undef AXI_R1_BEA_S6
`endif 

`ifdef AXI_R1_BSA_S7
  `undef AXI_R1_BSA_S7
`endif 

`ifdef AXI_R1_BEA_S7
  `undef AXI_R1_BEA_S7
`endif 

`ifdef AXI_R1_BSA_S8
  `undef AXI_R1_BSA_S8
`endif 

`ifdef AXI_R1_BEA_S8
  `undef AXI_R1_BEA_S8
`endif 

`ifdef AXI_R1_BSA_S9
  `undef AXI_R1_BSA_S9
`endif 

`ifdef AXI_R1_BEA_S9
  `undef AXI_R1_BEA_S9
`endif 

`ifdef AXI_R1_BSA_S10
  `undef AXI_R1_BSA_S10
`endif 

`ifdef AXI_R1_BEA_S10
  `undef AXI_R1_BEA_S10
`endif 

`ifdef AXI_R1_BSA_S11
  `undef AXI_R1_BSA_S11
`endif 

`ifdef AXI_R1_BEA_S11
  `undef AXI_R1_BEA_S11
`endif 

`ifdef AXI_R1_BSA_S12
  `undef AXI_R1_BSA_S12
`endif 

`ifdef AXI_R1_BEA_S12
  `undef AXI_R1_BEA_S12
`endif 

`ifdef AXI_R1_BSA_S13
  `undef AXI_R1_BSA_S13
`endif 

`ifdef AXI_R1_BEA_S13
  `undef AXI_R1_BEA_S13
`endif 

`ifdef AXI_R1_BSA_S14
  `undef AXI_R1_BSA_S14
`endif 

`ifdef AXI_R1_BEA_S14
  `undef AXI_R1_BEA_S14
`endif 

`ifdef AXI_R1_BSA_S15
  `undef AXI_R1_BSA_S15
`endif 

`ifdef AXI_R1_BEA_S15
  `undef AXI_R1_BEA_S15
`endif 

`ifdef AXI_R1_BSA_S16
  `undef AXI_R1_BSA_S16
`endif 

`ifdef AXI_R1_BEA_S16
  `undef AXI_R1_BEA_S16
`endif 

`ifdef AXI_R2_BSA_S1
  `undef AXI_R2_BSA_S1
`endif 

`ifdef AXI_R2_BEA_S1
  `undef AXI_R2_BEA_S1
`endif 

`ifdef AXI_R2_BSA_S2
  `undef AXI_R2_BSA_S2
`endif 

`ifdef AXI_R2_BEA_S2
  `undef AXI_R2_BEA_S2
`endif 

`ifdef AXI_R2_BSA_S3
  `undef AXI_R2_BSA_S3
`endif 

`ifdef AXI_R2_BEA_S3
  `undef AXI_R2_BEA_S3
`endif 

`ifdef AXI_R2_BSA_S4
  `undef AXI_R2_BSA_S4
`endif 

`ifdef AXI_R2_BEA_S4
  `undef AXI_R2_BEA_S4
`endif 

`ifdef AXI_R2_BSA_S5
  `undef AXI_R2_BSA_S5
`endif 

`ifdef AXI_R2_BEA_S5
  `undef AXI_R2_BEA_S5
`endif 

`ifdef AXI_R2_BSA_S6
  `undef AXI_R2_BSA_S6
`endif 

`ifdef AXI_R2_BEA_S6
  `undef AXI_R2_BEA_S6
`endif 

`ifdef AXI_R2_BSA_S7
  `undef AXI_R2_BSA_S7
`endif 

`ifdef AXI_R2_BEA_S7
  `undef AXI_R2_BEA_S7
`endif 

`ifdef AXI_R2_BSA_S8
  `undef AXI_R2_BSA_S8
`endif 

`ifdef AXI_R2_BEA_S8
  `undef AXI_R2_BEA_S8
`endif 

`ifdef AXI_R2_BSA_S9
  `undef AXI_R2_BSA_S9
`endif 

`ifdef AXI_R2_BEA_S9
  `undef AXI_R2_BEA_S9
`endif 

`ifdef AXI_R2_BSA_S10
  `undef AXI_R2_BSA_S10
`endif 

`ifdef AXI_R2_BEA_S10
  `undef AXI_R2_BEA_S10
`endif 

`ifdef AXI_R2_BSA_S11
  `undef AXI_R2_BSA_S11
`endif 

`ifdef AXI_R2_BEA_S11
  `undef AXI_R2_BEA_S11
`endif 

`ifdef AXI_R2_BSA_S12
  `undef AXI_R2_BSA_S12
`endif 

`ifdef AXI_R2_BEA_S12
  `undef AXI_R2_BEA_S12
`endif 

`ifdef AXI_R2_BSA_S13
  `undef AXI_R2_BSA_S13
`endif 

`ifdef AXI_R2_BEA_S13
  `undef AXI_R2_BEA_S13
`endif 

`ifdef AXI_R2_BSA_S14
  `undef AXI_R2_BSA_S14
`endif 

`ifdef AXI_R2_BEA_S14
  `undef AXI_R2_BEA_S14
`endif 

`ifdef AXI_R2_BSA_S15
  `undef AXI_R2_BSA_S15
`endif 

`ifdef AXI_R2_BEA_S15
  `undef AXI_R2_BEA_S15
`endif 

`ifdef AXI_R2_BSA_S16
  `undef AXI_R2_BSA_S16
`endif 

`ifdef AXI_R2_BEA_S16
  `undef AXI_R2_BEA_S16
`endif 

`ifdef AXI_R3_BSA_S1
  `undef AXI_R3_BSA_S1
`endif 

`ifdef AXI_R3_BEA_S1
  `undef AXI_R3_BEA_S1
`endif 

`ifdef AXI_R3_BSA_S2
  `undef AXI_R3_BSA_S2
`endif 

`ifdef AXI_R3_BEA_S2
  `undef AXI_R3_BEA_S2
`endif 

`ifdef AXI_R3_BSA_S3
  `undef AXI_R3_BSA_S3
`endif 

`ifdef AXI_R3_BEA_S3
  `undef AXI_R3_BEA_S3
`endif 

`ifdef AXI_R3_BSA_S4
  `undef AXI_R3_BSA_S4
`endif 

`ifdef AXI_R3_BEA_S4
  `undef AXI_R3_BEA_S4
`endif 

`ifdef AXI_R3_BSA_S5
  `undef AXI_R3_BSA_S5
`endif 

`ifdef AXI_R3_BEA_S5
  `undef AXI_R3_BEA_S5
`endif 

`ifdef AXI_R3_BSA_S6
  `undef AXI_R3_BSA_S6
`endif 

`ifdef AXI_R3_BEA_S6
  `undef AXI_R3_BEA_S6
`endif 

`ifdef AXI_R3_BSA_S7
  `undef AXI_R3_BSA_S7
`endif 

`ifdef AXI_R3_BEA_S7
  `undef AXI_R3_BEA_S7
`endif 

`ifdef AXI_R3_BSA_S8
  `undef AXI_R3_BSA_S8
`endif 

`ifdef AXI_R3_BEA_S8
  `undef AXI_R3_BEA_S8
`endif 

`ifdef AXI_R3_BSA_S9
  `undef AXI_R3_BSA_S9
`endif 

`ifdef AXI_R3_BEA_S9
  `undef AXI_R3_BEA_S9
`endif 

`ifdef AXI_R3_BSA_S10
  `undef AXI_R3_BSA_S10
`endif 

`ifdef AXI_R3_BEA_S10
  `undef AXI_R3_BEA_S10
`endif 

`ifdef AXI_R3_BSA_S11
  `undef AXI_R3_BSA_S11
`endif 

`ifdef AXI_R3_BEA_S11
  `undef AXI_R3_BEA_S11
`endif 

`ifdef AXI_R3_BSA_S12
  `undef AXI_R3_BSA_S12
`endif 

`ifdef AXI_R3_BEA_S12
  `undef AXI_R3_BEA_S12
`endif 

`ifdef AXI_R3_BSA_S13
  `undef AXI_R3_BSA_S13
`endif 

`ifdef AXI_R3_BEA_S13
  `undef AXI_R3_BEA_S13
`endif 

`ifdef AXI_R3_BSA_S14
  `undef AXI_R3_BSA_S14
`endif 

`ifdef AXI_R3_BEA_S14
  `undef AXI_R3_BEA_S14
`endif 

`ifdef AXI_R3_BSA_S15
  `undef AXI_R3_BSA_S15
`endif 

`ifdef AXI_R3_BEA_S15
  `undef AXI_R3_BEA_S15
`endif 

`ifdef AXI_R3_BSA_S16
  `undef AXI_R3_BSA_S16
`endif 

`ifdef AXI_R3_BEA_S16
  `undef AXI_R3_BEA_S16
`endif 

`ifdef AXI_R4_BSA_S1
  `undef AXI_R4_BSA_S1
`endif 

`ifdef AXI_R4_BEA_S1
  `undef AXI_R4_BEA_S1
`endif 

`ifdef AXI_R4_BSA_S2
  `undef AXI_R4_BSA_S2
`endif 

`ifdef AXI_R4_BEA_S2
  `undef AXI_R4_BEA_S2
`endif 

`ifdef AXI_R4_BSA_S3
  `undef AXI_R4_BSA_S3
`endif 

`ifdef AXI_R4_BEA_S3
  `undef AXI_R4_BEA_S3
`endif 

`ifdef AXI_R4_BSA_S4
  `undef AXI_R4_BSA_S4
`endif 

`ifdef AXI_R4_BEA_S4
  `undef AXI_R4_BEA_S4
`endif 

`ifdef AXI_R4_BSA_S5
  `undef AXI_R4_BSA_S5
`endif 

`ifdef AXI_R4_BEA_S5
  `undef AXI_R4_BEA_S5
`endif 

`ifdef AXI_R4_BSA_S6
  `undef AXI_R4_BSA_S6
`endif 

`ifdef AXI_R4_BEA_S6
  `undef AXI_R4_BEA_S6
`endif 

`ifdef AXI_R4_BSA_S7
  `undef AXI_R4_BSA_S7
`endif 

`ifdef AXI_R4_BEA_S7
  `undef AXI_R4_BEA_S7
`endif 

`ifdef AXI_R4_BSA_S8
  `undef AXI_R4_BSA_S8
`endif 

`ifdef AXI_R4_BEA_S8
  `undef AXI_R4_BEA_S8
`endif 

`ifdef AXI_R4_BSA_S9
  `undef AXI_R4_BSA_S9
`endif 

`ifdef AXI_R4_BEA_S9
  `undef AXI_R4_BEA_S9
`endif 

`ifdef AXI_R4_BSA_S10
  `undef AXI_R4_BSA_S10
`endif 

`ifdef AXI_R4_BEA_S10
  `undef AXI_R4_BEA_S10
`endif 

`ifdef AXI_R4_BSA_S11
  `undef AXI_R4_BSA_S11
`endif 

`ifdef AXI_R4_BEA_S11
  `undef AXI_R4_BEA_S11
`endif 

`ifdef AXI_R4_BSA_S12
  `undef AXI_R4_BSA_S12
`endif 

`ifdef AXI_R4_BEA_S12
  `undef AXI_R4_BEA_S12
`endif 

`ifdef AXI_R4_BSA_S13
  `undef AXI_R4_BSA_S13
`endif 

`ifdef AXI_R4_BEA_S13
  `undef AXI_R4_BEA_S13
`endif 

`ifdef AXI_R4_BSA_S14
  `undef AXI_R4_BSA_S14
`endif 

`ifdef AXI_R4_BEA_S14
  `undef AXI_R4_BEA_S14
`endif 

`ifdef AXI_R4_BSA_S15
  `undef AXI_R4_BSA_S15
`endif 

`ifdef AXI_R4_BEA_S15
  `undef AXI_R4_BEA_S15
`endif 

`ifdef AXI_R4_BSA_S16
  `undef AXI_R4_BSA_S16
`endif 

`ifdef AXI_R4_BEA_S16
  `undef AXI_R4_BEA_S16
`endif 

`ifdef AXI_R5_BSA_S1
  `undef AXI_R5_BSA_S1
`endif 

`ifdef AXI_R5_BEA_S1
  `undef AXI_R5_BEA_S1
`endif 

`ifdef AXI_R5_BSA_S2
  `undef AXI_R5_BSA_S2
`endif 

`ifdef AXI_R5_BEA_S2
  `undef AXI_R5_BEA_S2
`endif 

`ifdef AXI_R5_BSA_S3
  `undef AXI_R5_BSA_S3
`endif 

`ifdef AXI_R5_BEA_S3
  `undef AXI_R5_BEA_S3
`endif 

`ifdef AXI_R5_BSA_S4
  `undef AXI_R5_BSA_S4
`endif 

`ifdef AXI_R5_BEA_S4
  `undef AXI_R5_BEA_S4
`endif 

`ifdef AXI_R5_BSA_S5
  `undef AXI_R5_BSA_S5
`endif 

`ifdef AXI_R5_BEA_S5
  `undef AXI_R5_BEA_S5
`endif 

`ifdef AXI_R5_BSA_S6
  `undef AXI_R5_BSA_S6
`endif 

`ifdef AXI_R5_BEA_S6
  `undef AXI_R5_BEA_S6
`endif 

`ifdef AXI_R5_BSA_S7
  `undef AXI_R5_BSA_S7
`endif 

`ifdef AXI_R5_BEA_S7
  `undef AXI_R5_BEA_S7
`endif 

`ifdef AXI_R5_BSA_S8
  `undef AXI_R5_BSA_S8
`endif 

`ifdef AXI_R5_BEA_S8
  `undef AXI_R5_BEA_S8
`endif 

`ifdef AXI_R5_BSA_S9
  `undef AXI_R5_BSA_S9
`endif 

`ifdef AXI_R5_BEA_S9
  `undef AXI_R5_BEA_S9
`endif 

`ifdef AXI_R5_BSA_S10
  `undef AXI_R5_BSA_S10
`endif 

`ifdef AXI_R5_BEA_S10
  `undef AXI_R5_BEA_S10
`endif 

`ifdef AXI_R5_BSA_S11
  `undef AXI_R5_BSA_S11
`endif 

`ifdef AXI_R5_BEA_S11
  `undef AXI_R5_BEA_S11
`endif 

`ifdef AXI_R5_BSA_S12
  `undef AXI_R5_BSA_S12
`endif 

`ifdef AXI_R5_BEA_S12
  `undef AXI_R5_BEA_S12
`endif 

`ifdef AXI_R5_BSA_S13
  `undef AXI_R5_BSA_S13
`endif 

`ifdef AXI_R5_BEA_S13
  `undef AXI_R5_BEA_S13
`endif 

`ifdef AXI_R5_BSA_S14
  `undef AXI_R5_BSA_S14
`endif 

`ifdef AXI_R5_BEA_S14
  `undef AXI_R5_BEA_S14
`endif 

`ifdef AXI_R5_BSA_S15
  `undef AXI_R5_BSA_S15
`endif 

`ifdef AXI_R5_BEA_S15
  `undef AXI_R5_BEA_S15
`endif 

`ifdef AXI_R5_BSA_S16
  `undef AXI_R5_BSA_S16
`endif 

`ifdef AXI_R5_BEA_S16
  `undef AXI_R5_BEA_S16
`endif 

`ifdef AXI_R6_BSA_S1
  `undef AXI_R6_BSA_S1
`endif 

`ifdef AXI_R6_BEA_S1
  `undef AXI_R6_BEA_S1
`endif 

`ifdef AXI_R6_BSA_S2
  `undef AXI_R6_BSA_S2
`endif 

`ifdef AXI_R6_BEA_S2
  `undef AXI_R6_BEA_S2
`endif 

`ifdef AXI_R6_BSA_S3
  `undef AXI_R6_BSA_S3
`endif 

`ifdef AXI_R6_BEA_S3
  `undef AXI_R6_BEA_S3
`endif 

`ifdef AXI_R6_BSA_S4
  `undef AXI_R6_BSA_S4
`endif 

`ifdef AXI_R6_BEA_S4
  `undef AXI_R6_BEA_S4
`endif 

`ifdef AXI_R6_BSA_S5
  `undef AXI_R6_BSA_S5
`endif 

`ifdef AXI_R6_BEA_S5
  `undef AXI_R6_BEA_S5
`endif 

`ifdef AXI_R6_BSA_S6
  `undef AXI_R6_BSA_S6
`endif 

`ifdef AXI_R6_BEA_S6
  `undef AXI_R6_BEA_S6
`endif 

`ifdef AXI_R6_BSA_S7
  `undef AXI_R6_BSA_S7
`endif 

`ifdef AXI_R6_BEA_S7
  `undef AXI_R6_BEA_S7
`endif 

`ifdef AXI_R6_BSA_S8
  `undef AXI_R6_BSA_S8
`endif 

`ifdef AXI_R6_BEA_S8
  `undef AXI_R6_BEA_S8
`endif 

`ifdef AXI_R6_BSA_S9
  `undef AXI_R6_BSA_S9
`endif 

`ifdef AXI_R6_BEA_S9
  `undef AXI_R6_BEA_S9
`endif 

`ifdef AXI_R6_BSA_S10
  `undef AXI_R6_BSA_S10
`endif 

`ifdef AXI_R6_BEA_S10
  `undef AXI_R6_BEA_S10
`endif 

`ifdef AXI_R6_BSA_S11
  `undef AXI_R6_BSA_S11
`endif 

`ifdef AXI_R6_BEA_S11
  `undef AXI_R6_BEA_S11
`endif 

`ifdef AXI_R6_BSA_S12
  `undef AXI_R6_BSA_S12
`endif 

`ifdef AXI_R6_BEA_S12
  `undef AXI_R6_BEA_S12
`endif 

`ifdef AXI_R6_BSA_S13
  `undef AXI_R6_BSA_S13
`endif 

`ifdef AXI_R6_BEA_S13
  `undef AXI_R6_BEA_S13
`endif 

`ifdef AXI_R6_BSA_S14
  `undef AXI_R6_BSA_S14
`endif 

`ifdef AXI_R6_BEA_S14
  `undef AXI_R6_BEA_S14
`endif 

`ifdef AXI_R6_BSA_S15
  `undef AXI_R6_BSA_S15
`endif 

`ifdef AXI_R6_BEA_S15
  `undef AXI_R6_BEA_S15
`endif 

`ifdef AXI_R6_BSA_S16
  `undef AXI_R6_BSA_S16
`endif 

`ifdef AXI_R6_BEA_S16
  `undef AXI_R6_BEA_S16
`endif 

`ifdef AXI_R7_BSA_S1
  `undef AXI_R7_BSA_S1
`endif 

`ifdef AXI_R7_BEA_S1
  `undef AXI_R7_BEA_S1
`endif 

`ifdef AXI_R7_BSA_S2
  `undef AXI_R7_BSA_S2
`endif 

`ifdef AXI_R7_BEA_S2
  `undef AXI_R7_BEA_S2
`endif 

`ifdef AXI_R7_BSA_S3
  `undef AXI_R7_BSA_S3
`endif 

`ifdef AXI_R7_BEA_S3
  `undef AXI_R7_BEA_S3
`endif 

`ifdef AXI_R7_BSA_S4
  `undef AXI_R7_BSA_S4
`endif 

`ifdef AXI_R7_BEA_S4
  `undef AXI_R7_BEA_S4
`endif 

`ifdef AXI_R7_BSA_S5
  `undef AXI_R7_BSA_S5
`endif 

`ifdef AXI_R7_BEA_S5
  `undef AXI_R7_BEA_S5
`endif 

`ifdef AXI_R7_BSA_S6
  `undef AXI_R7_BSA_S6
`endif 

`ifdef AXI_R7_BEA_S6
  `undef AXI_R7_BEA_S6
`endif 

`ifdef AXI_R7_BSA_S7
  `undef AXI_R7_BSA_S7
`endif 

`ifdef AXI_R7_BEA_S7
  `undef AXI_R7_BEA_S7
`endif 

`ifdef AXI_R7_BSA_S8
  `undef AXI_R7_BSA_S8
`endif 

`ifdef AXI_R7_BEA_S8
  `undef AXI_R7_BEA_S8
`endif 

`ifdef AXI_R7_BSA_S9
  `undef AXI_R7_BSA_S9
`endif 

`ifdef AXI_R7_BEA_S9
  `undef AXI_R7_BEA_S9
`endif 

`ifdef AXI_R7_BSA_S10
  `undef AXI_R7_BSA_S10
`endif 

`ifdef AXI_R7_BEA_S10
  `undef AXI_R7_BEA_S10
`endif 

`ifdef AXI_R7_BSA_S11
  `undef AXI_R7_BSA_S11
`endif 

`ifdef AXI_R7_BEA_S11
  `undef AXI_R7_BEA_S11
`endif 

`ifdef AXI_R7_BSA_S12
  `undef AXI_R7_BSA_S12
`endif 

`ifdef AXI_R7_BEA_S12
  `undef AXI_R7_BEA_S12
`endif 

`ifdef AXI_R7_BSA_S13
  `undef AXI_R7_BSA_S13
`endif 

`ifdef AXI_R7_BEA_S13
  `undef AXI_R7_BEA_S13
`endif 

`ifdef AXI_R7_BSA_S14
  `undef AXI_R7_BSA_S14
`endif 

`ifdef AXI_R7_BEA_S14
  `undef AXI_R7_BEA_S14
`endif 

`ifdef AXI_R7_BSA_S15
  `undef AXI_R7_BSA_S15
`endif 

`ifdef AXI_R7_BEA_S15
  `undef AXI_R7_BEA_S15
`endif 

`ifdef AXI_R7_BSA_S16
  `undef AXI_R7_BSA_S16
`endif 

`ifdef AXI_R7_BEA_S16
  `undef AXI_R7_BEA_S16
`endif 

`ifdef AXI_R8_BSA_S1
  `undef AXI_R8_BSA_S1
`endif 

`ifdef AXI_R8_BEA_S1
  `undef AXI_R8_BEA_S1
`endif 

`ifdef AXI_R8_BSA_S2
  `undef AXI_R8_BSA_S2
`endif 

`ifdef AXI_R8_BEA_S2
  `undef AXI_R8_BEA_S2
`endif 

`ifdef AXI_R8_BSA_S3
  `undef AXI_R8_BSA_S3
`endif 

`ifdef AXI_R8_BEA_S3
  `undef AXI_R8_BEA_S3
`endif 

`ifdef AXI_R8_BSA_S4
  `undef AXI_R8_BSA_S4
`endif 

`ifdef AXI_R8_BEA_S4
  `undef AXI_R8_BEA_S4
`endif 

`ifdef AXI_R8_BSA_S5
  `undef AXI_R8_BSA_S5
`endif 

`ifdef AXI_R8_BEA_S5
  `undef AXI_R8_BEA_S5
`endif 

`ifdef AXI_R8_BSA_S6
  `undef AXI_R8_BSA_S6
`endif 

`ifdef AXI_R8_BEA_S6
  `undef AXI_R8_BEA_S6
`endif 

`ifdef AXI_R8_BSA_S7
  `undef AXI_R8_BSA_S7
`endif 

`ifdef AXI_R8_BEA_S7
  `undef AXI_R8_BEA_S7
`endif 

`ifdef AXI_R8_BSA_S8
  `undef AXI_R8_BSA_S8
`endif 

`ifdef AXI_R8_BEA_S8
  `undef AXI_R8_BEA_S8
`endif 

`ifdef AXI_R8_BSA_S9
  `undef AXI_R8_BSA_S9
`endif 

`ifdef AXI_R8_BEA_S9
  `undef AXI_R8_BEA_S9
`endif 

`ifdef AXI_R8_BSA_S10
  `undef AXI_R8_BSA_S10
`endif 

`ifdef AXI_R8_BEA_S10
  `undef AXI_R8_BEA_S10
`endif 

`ifdef AXI_R8_BSA_S11
  `undef AXI_R8_BSA_S11
`endif 

`ifdef AXI_R8_BEA_S11
  `undef AXI_R8_BEA_S11
`endif 

`ifdef AXI_R8_BSA_S12
  `undef AXI_R8_BSA_S12
`endif 

`ifdef AXI_R8_BEA_S12
  `undef AXI_R8_BEA_S12
`endif 

`ifdef AXI_R8_BSA_S13
  `undef AXI_R8_BSA_S13
`endif 

`ifdef AXI_R8_BEA_S13
  `undef AXI_R8_BEA_S13
`endif 

`ifdef AXI_R8_BSA_S14
  `undef AXI_R8_BSA_S14
`endif 

`ifdef AXI_R8_BEA_S14
  `undef AXI_R8_BEA_S14
`endif 

`ifdef AXI_R8_BSA_S15
  `undef AXI_R8_BSA_S15
`endif 

`ifdef AXI_R8_BEA_S15
  `undef AXI_R8_BEA_S15
`endif 

`ifdef AXI_R8_BSA_S16
  `undef AXI_R8_BSA_S16
`endif 

`ifdef AXI_R8_BEA_S16
  `undef AXI_R8_BEA_S16
`endif 

`ifdef AXI_AR_PYLD_M_W
  `undef AXI_AR_PYLD_M_W
`endif 

`ifdef AXI_AW_PYLD_M_W
  `undef AXI_AW_PYLD_M_W
`endif 

`ifdef AXI_W_PYLD_M_W
  `undef AXI_W_PYLD_M_W
`endif 

`ifdef AXI_R_PYLD_M_W
  `undef AXI_R_PYLD_M_W
`endif 

`ifdef AXI_B_PYLD_M_W
  `undef AXI_B_PYLD_M_W
`endif 

`ifdef AXI_AR_PYLD_S_W
  `undef AXI_AR_PYLD_S_W
`endif 

`ifdef AXI_AW_PYLD_S_W
  `undef AXI_AW_PYLD_S_W
`endif 

`ifdef AXI_W_PYLD_S_W
  `undef AXI_W_PYLD_S_W
`endif 

`ifdef AXI_R_PYLD_S_W
  `undef AXI_R_PYLD_S_W
`endif 

`ifdef AXI_B_PYLD_S_W
  `undef AXI_B_PYLD_S_W
`endif 

`ifdef AXI_HAS_S0
  `undef AXI_HAS_S0
`endif 

`ifdef AXI_HAS_S1
  `undef AXI_HAS_S1
`endif 

`ifdef AXI_HAS_S2
  `undef AXI_HAS_S2
`endif 

`ifdef AXI_HAS_S3
  `undef AXI_HAS_S3
`endif 

`ifdef AXI_HAS_M1
  `undef AXI_HAS_M1
`endif 

`ifdef AXI_HAS_M2
  `undef AXI_HAS_M2
`endif 

`ifdef AXI_NMV_S0
  `undef AXI_NMV_S0
`endif 

`ifdef AXI_SYS_NUM_FOR_M1
  `undef AXI_SYS_NUM_FOR_M1
`endif 

`ifdef AXI_SYS_NUM_FOR_M2
  `undef AXI_SYS_NUM_FOR_M2
`endif 

`ifdef AXI_SYS_NUM_FOR_M3
  `undef AXI_SYS_NUM_FOR_M3
`endif 

`ifdef AXI_SYS_NUM_FOR_M4
  `undef AXI_SYS_NUM_FOR_M4
`endif 

`ifdef AXI_SYS_NUM_FOR_M5
  `undef AXI_SYS_NUM_FOR_M5
`endif 

`ifdef AXI_SYS_NUM_FOR_M6
  `undef AXI_SYS_NUM_FOR_M6
`endif 

`ifdef AXI_SYS_NUM_FOR_M7
  `undef AXI_SYS_NUM_FOR_M7
`endif 

`ifdef AXI_SYS_NUM_FOR_M8
  `undef AXI_SYS_NUM_FOR_M8
`endif 

`ifdef AXI_SYS_NUM_FOR_M9
  `undef AXI_SYS_NUM_FOR_M9
`endif 

`ifdef AXI_SYS_NUM_FOR_M10
  `undef AXI_SYS_NUM_FOR_M10
`endif 

`ifdef AXI_SYS_NUM_FOR_M11
  `undef AXI_SYS_NUM_FOR_M11
`endif 

`ifdef AXI_SYS_NUM_FOR_M12
  `undef AXI_SYS_NUM_FOR_M12
`endif 

`ifdef AXI_SYS_NUM_FOR_M13
  `undef AXI_SYS_NUM_FOR_M13
`endif 

`ifdef AXI_SYS_NUM_FOR_M14
  `undef AXI_SYS_NUM_FOR_M14
`endif 

`ifdef AXI_SYS_NUM_FOR_M15
  `undef AXI_SYS_NUM_FOR_M15
`endif 

`ifdef AXI_SYS_NUM_FOR_M16
  `undef AXI_SYS_NUM_FOR_M16
`endif 

`ifdef AXI_NUM_ICM
  `undef AXI_NUM_ICM
`endif 

`ifdef AXI_ACC_NON_LCL_SLV_S1
  `undef AXI_ACC_NON_LCL_SLV_S1
`endif 

`ifdef AXI_ACC_NON_LCL_SLV_S2
  `undef AXI_ACC_NON_LCL_SLV_S2
`endif 

`ifdef AXI_ACC_NON_LCL_SLV_S3
  `undef AXI_ACC_NON_LCL_SLV_S3
`endif 

`ifdef AXI_ACC_NON_LCL_SLV_S4
  `undef AXI_ACC_NON_LCL_SLV_S4
`endif 

`ifdef AXI_ACC_NON_LCL_SLV_S5
  `undef AXI_ACC_NON_LCL_SLV_S5
`endif 

`ifdef AXI_ACC_NON_LCL_SLV_S6
  `undef AXI_ACC_NON_LCL_SLV_S6
`endif 

`ifdef AXI_ACC_NON_LCL_SLV_S7
  `undef AXI_ACC_NON_LCL_SLV_S7
`endif 

`ifdef AXI_ACC_NON_LCL_SLV_S8
  `undef AXI_ACC_NON_LCL_SLV_S8
`endif 

`ifdef AXI_ACC_NON_LCL_SLV_S9
  `undef AXI_ACC_NON_LCL_SLV_S9
`endif 

`ifdef AXI_ACC_NON_LCL_SLV_S10
  `undef AXI_ACC_NON_LCL_SLV_S10
`endif 

`ifdef AXI_ACC_NON_LCL_SLV_S11
  `undef AXI_ACC_NON_LCL_SLV_S11
`endif 

`ifdef AXI_ACC_NON_LCL_SLV_S12
  `undef AXI_ACC_NON_LCL_SLV_S12
`endif 

`ifdef AXI_ACC_NON_LCL_SLV_S13
  `undef AXI_ACC_NON_LCL_SLV_S13
`endif 

`ifdef AXI_ACC_NON_LCL_SLV_S14
  `undef AXI_ACC_NON_LCL_SLV_S14
`endif 

`ifdef AXI_ACC_NON_LCL_SLV_S15
  `undef AXI_ACC_NON_LCL_SLV_S15
`endif 

`ifdef AXI_ACC_NON_LCL_SLV_S16
  `undef AXI_ACC_NON_LCL_SLV_S16
`endif 

`ifdef AXI_IS_ICM_M1
  `undef AXI_IS_ICM_M1
`endif 

`ifdef AXI_IS_ICM_M2
  `undef AXI_IS_ICM_M2
`endif 

`ifdef AXI_IS_ICM_M3
  `undef AXI_IS_ICM_M3
`endif 

`ifdef AXI_IS_ICM_M4
  `undef AXI_IS_ICM_M4
`endif 

`ifdef AXI_IS_ICM_M5
  `undef AXI_IS_ICM_M5
`endif 

`ifdef AXI_IS_ICM_M6
  `undef AXI_IS_ICM_M6
`endif 

`ifdef AXI_IS_ICM_M7
  `undef AXI_IS_ICM_M7
`endif 

`ifdef AXI_IS_ICM_M8
  `undef AXI_IS_ICM_M8
`endif 

`ifdef AXI_IS_ICM_M9
  `undef AXI_IS_ICM_M9
`endif 

`ifdef AXI_IS_ICM_M10
  `undef AXI_IS_ICM_M10
`endif 

`ifdef AXI_IS_ICM_M11
  `undef AXI_IS_ICM_M11
`endif 

`ifdef AXI_IS_ICM_M12
  `undef AXI_IS_ICM_M12
`endif 

`ifdef AXI_IS_ICM_M13
  `undef AXI_IS_ICM_M13
`endif 

`ifdef AXI_IS_ICM_M14
  `undef AXI_IS_ICM_M14
`endif 

`ifdef AXI_IS_ICM_M15
  `undef AXI_IS_ICM_M15
`endif 

`ifdef AXI_IS_ICM_M16
  `undef AXI_IS_ICM_M16
`endif 

`ifdef AXI_HAS_ICM1
  `undef AXI_HAS_ICM1
`endif 

`ifdef AXI_HAS_ICM2
  `undef AXI_HAS_ICM2
`endif 

`ifdef AXI_HAS_ICM3
  `undef AXI_HAS_ICM3
`endif 

`ifdef AXI_HAS_ICM4
  `undef AXI_HAS_ICM4
`endif 

`ifdef AXI_IDW_M1
  `undef AXI_IDW_M1
`endif 

`ifdef AXI_IDW_M2
  `undef AXI_IDW_M2
`endif 

`ifdef AXI_IDW_M3
  `undef AXI_IDW_M3
`endif 

`ifdef AXI_IDW_M4
  `undef AXI_IDW_M4
`endif 

`ifdef AXI_NUM_MST_THRU_ICM1
  `undef AXI_NUM_MST_THRU_ICM1
`endif 

`ifdef AXI_NUM_MST_THRU_ICM2
  `undef AXI_NUM_MST_THRU_ICM2
`endif 

`ifdef AXI_NUM_MST_THRU_ICM3
  `undef AXI_NUM_MST_THRU_ICM3
`endif 

`ifdef AXI_NUM_MST_THRU_ICM4
  `undef AXI_NUM_MST_THRU_ICM4
`endif 

`ifdef AXI_ALLOW_MST1_ICM1
  `undef AXI_ALLOW_MST1_ICM1
`endif 

`ifdef AXI_ALLOW_MST2_ICM1
  `undef AXI_ALLOW_MST2_ICM1
`endif 

`ifdef AXI_ALLOW_MST3_ICM1
  `undef AXI_ALLOW_MST3_ICM1
`endif 

`ifdef AXI_ALLOW_MST4_ICM1
  `undef AXI_ALLOW_MST4_ICM1
`endif 

`ifdef AXI_ALLOW_MST5_ICM1
  `undef AXI_ALLOW_MST5_ICM1
`endif 

`ifdef AXI_ALLOW_MST6_ICM1
  `undef AXI_ALLOW_MST6_ICM1
`endif 

`ifdef AXI_ALLOW_MST7_ICM1
  `undef AXI_ALLOW_MST7_ICM1
`endif 

`ifdef AXI_ALLOW_MST8_ICM1
  `undef AXI_ALLOW_MST8_ICM1
`endif 

`ifdef AXI_ALLOW_MST1_ICM2
  `undef AXI_ALLOW_MST1_ICM2
`endif 

`ifdef AXI_ALLOW_MST2_ICM2
  `undef AXI_ALLOW_MST2_ICM2
`endif 

`ifdef AXI_ALLOW_MST3_ICM2
  `undef AXI_ALLOW_MST3_ICM2
`endif 

`ifdef AXI_ALLOW_MST4_ICM2
  `undef AXI_ALLOW_MST4_ICM2
`endif 

`ifdef AXI_ALLOW_MST5_ICM2
  `undef AXI_ALLOW_MST5_ICM2
`endif 

`ifdef AXI_ALLOW_MST6_ICM2
  `undef AXI_ALLOW_MST6_ICM2
`endif 

`ifdef AXI_ALLOW_MST7_ICM2
  `undef AXI_ALLOW_MST7_ICM2
`endif 

`ifdef AXI_ALLOW_MST8_ICM2
  `undef AXI_ALLOW_MST8_ICM2
`endif 

`ifdef AXI_ALLOW_MST1_ICM3
  `undef AXI_ALLOW_MST1_ICM3
`endif 

`ifdef AXI_ALLOW_MST2_ICM3
  `undef AXI_ALLOW_MST2_ICM3
`endif 

`ifdef AXI_ALLOW_MST3_ICM3
  `undef AXI_ALLOW_MST3_ICM3
`endif 

`ifdef AXI_ALLOW_MST4_ICM3
  `undef AXI_ALLOW_MST4_ICM3
`endif 

`ifdef AXI_ALLOW_MST5_ICM3
  `undef AXI_ALLOW_MST5_ICM3
`endif 

`ifdef AXI_ALLOW_MST6_ICM3
  `undef AXI_ALLOW_MST6_ICM3
`endif 

`ifdef AXI_ALLOW_MST7_ICM3
  `undef AXI_ALLOW_MST7_ICM3
`endif 

`ifdef AXI_ALLOW_MST8_ICM3
  `undef AXI_ALLOW_MST8_ICM3
`endif 

`ifdef AXI_ALLOW_MST1_ICM4
  `undef AXI_ALLOW_MST1_ICM4
`endif 

`ifdef AXI_ALLOW_MST2_ICM4
  `undef AXI_ALLOW_MST2_ICM4
`endif 

`ifdef AXI_ALLOW_MST3_ICM4
  `undef AXI_ALLOW_MST3_ICM4
`endif 

`ifdef AXI_ALLOW_MST4_ICM4
  `undef AXI_ALLOW_MST4_ICM4
`endif 

`ifdef AXI_ALLOW_MST5_ICM4
  `undef AXI_ALLOW_MST5_ICM4
`endif 

`ifdef AXI_ALLOW_MST6_ICM4
  `undef AXI_ALLOW_MST6_ICM4
`endif 

`ifdef AXI_ALLOW_MST7_ICM4
  `undef AXI_ALLOW_MST7_ICM4
`endif 

`ifdef AXI_ALLOW_MST8_ICM4
  `undef AXI_ALLOW_MST8_ICM4
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M1
  `undef AXI_PNUM_FOR_SYS_NUM_M1
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M2
  `undef AXI_PNUM_FOR_SYS_NUM_M2
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M3
  `undef AXI_PNUM_FOR_SYS_NUM_M3
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M4
  `undef AXI_PNUM_FOR_SYS_NUM_M4
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M5
  `undef AXI_PNUM_FOR_SYS_NUM_M5
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M6
  `undef AXI_PNUM_FOR_SYS_NUM_M6
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M7
  `undef AXI_PNUM_FOR_SYS_NUM_M7
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M8
  `undef AXI_PNUM_FOR_SYS_NUM_M8
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M9
  `undef AXI_PNUM_FOR_SYS_NUM_M9
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M10
  `undef AXI_PNUM_FOR_SYS_NUM_M10
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M11
  `undef AXI_PNUM_FOR_SYS_NUM_M11
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M12
  `undef AXI_PNUM_FOR_SYS_NUM_M12
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M13
  `undef AXI_PNUM_FOR_SYS_NUM_M13
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M14
  `undef AXI_PNUM_FOR_SYS_NUM_M14
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M15
  `undef AXI_PNUM_FOR_SYS_NUM_M15
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M16
  `undef AXI_PNUM_FOR_SYS_NUM_M16
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M17
  `undef AXI_PNUM_FOR_SYS_NUM_M17
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M18
  `undef AXI_PNUM_FOR_SYS_NUM_M18
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M19
  `undef AXI_PNUM_FOR_SYS_NUM_M19
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M20
  `undef AXI_PNUM_FOR_SYS_NUM_M20
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M21
  `undef AXI_PNUM_FOR_SYS_NUM_M21
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M22
  `undef AXI_PNUM_FOR_SYS_NUM_M22
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M23
  `undef AXI_PNUM_FOR_SYS_NUM_M23
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M24
  `undef AXI_PNUM_FOR_SYS_NUM_M24
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M25
  `undef AXI_PNUM_FOR_SYS_NUM_M25
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M26
  `undef AXI_PNUM_FOR_SYS_NUM_M26
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M27
  `undef AXI_PNUM_FOR_SYS_NUM_M27
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M28
  `undef AXI_PNUM_FOR_SYS_NUM_M28
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M29
  `undef AXI_PNUM_FOR_SYS_NUM_M29
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M30
  `undef AXI_PNUM_FOR_SYS_NUM_M30
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M31
  `undef AXI_PNUM_FOR_SYS_NUM_M31
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M32
  `undef AXI_PNUM_FOR_SYS_NUM_M32
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M33
  `undef AXI_PNUM_FOR_SYS_NUM_M33
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M34
  `undef AXI_PNUM_FOR_SYS_NUM_M34
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M35
  `undef AXI_PNUM_FOR_SYS_NUM_M35
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M36
  `undef AXI_PNUM_FOR_SYS_NUM_M36
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M37
  `undef AXI_PNUM_FOR_SYS_NUM_M37
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M38
  `undef AXI_PNUM_FOR_SYS_NUM_M38
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M39
  `undef AXI_PNUM_FOR_SYS_NUM_M39
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M40
  `undef AXI_PNUM_FOR_SYS_NUM_M40
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M41
  `undef AXI_PNUM_FOR_SYS_NUM_M41
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M42
  `undef AXI_PNUM_FOR_SYS_NUM_M42
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M43
  `undef AXI_PNUM_FOR_SYS_NUM_M43
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M44
  `undef AXI_PNUM_FOR_SYS_NUM_M44
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M45
  `undef AXI_PNUM_FOR_SYS_NUM_M45
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M46
  `undef AXI_PNUM_FOR_SYS_NUM_M46
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M47
  `undef AXI_PNUM_FOR_SYS_NUM_M47
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M48
  `undef AXI_PNUM_FOR_SYS_NUM_M48
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M49
  `undef AXI_PNUM_FOR_SYS_NUM_M49
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M50
  `undef AXI_PNUM_FOR_SYS_NUM_M50
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M51
  `undef AXI_PNUM_FOR_SYS_NUM_M51
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M52
  `undef AXI_PNUM_FOR_SYS_NUM_M52
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M53
  `undef AXI_PNUM_FOR_SYS_NUM_M53
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M54
  `undef AXI_PNUM_FOR_SYS_NUM_M54
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M55
  `undef AXI_PNUM_FOR_SYS_NUM_M55
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M56
  `undef AXI_PNUM_FOR_SYS_NUM_M56
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M57
  `undef AXI_PNUM_FOR_SYS_NUM_M57
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M58
  `undef AXI_PNUM_FOR_SYS_NUM_M58
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M59
  `undef AXI_PNUM_FOR_SYS_NUM_M59
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M60
  `undef AXI_PNUM_FOR_SYS_NUM_M60
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M61
  `undef AXI_PNUM_FOR_SYS_NUM_M61
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M62
  `undef AXI_PNUM_FOR_SYS_NUM_M62
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M63
  `undef AXI_PNUM_FOR_SYS_NUM_M63
`endif 

`ifdef AXI_PNUM_FOR_SYS_NUM_M64
  `undef AXI_PNUM_FOR_SYS_NUM_M64
`endif 

`ifdef AXI_QOS
  `undef AXI_QOS
`endif 

`ifdef AXI_SRC_LICENSE_CHK
  `undef AXI_SRC_LICENSE_CHK
`endif 

`ifdef AXI_NSPV_M1_AR_QOSARB
  `undef AXI_NSPV_M1_AR_QOSARB
`endif 

`ifdef AXI_NSPV_M2_AR_QOSARB
  `undef AXI_NSPV_M2_AR_QOSARB
`endif 

`ifdef AXI_NSPV_M3_AR_QOSARB
  `undef AXI_NSPV_M3_AR_QOSARB
`endif 

`ifdef AXI_NSPV_M4_AR_QOSARB
  `undef AXI_NSPV_M4_AR_QOSARB
`endif 

`ifdef AXI_NSPV_M5_AR_QOSARB
  `undef AXI_NSPV_M5_AR_QOSARB
`endif 

`ifdef AXI_NSPV_M6_AR_QOSARB
  `undef AXI_NSPV_M6_AR_QOSARB
`endif 

`ifdef AXI_NSPV_M7_AR_QOSARB
  `undef AXI_NSPV_M7_AR_QOSARB
`endif 

`ifdef AXI_NSPV_M8_AR_QOSARB
  `undef AXI_NSPV_M8_AR_QOSARB
`endif 

`ifdef AXI_NSPV_M9_AR_QOSARB
  `undef AXI_NSPV_M9_AR_QOSARB
`endif 

`ifdef AXI_NSPV_M10_AR_QOSARB
  `undef AXI_NSPV_M10_AR_QOSARB
`endif 

`ifdef AXI_NSPV_M11_AR_QOSARB
  `undef AXI_NSPV_M11_AR_QOSARB
`endif 

`ifdef AXI_NSPV_M12_AR_QOSARB
  `undef AXI_NSPV_M12_AR_QOSARB
`endif 

`ifdef AXI_NSPV_M13_AR_QOSARB
  `undef AXI_NSPV_M13_AR_QOSARB
`endif 

`ifdef AXI_NSPV_M14_AR_QOSARB
  `undef AXI_NSPV_M14_AR_QOSARB
`endif 

`ifdef AXI_NSPV_M15_AR_QOSARB
  `undef AXI_NSPV_M15_AR_QOSARB
`endif 

`ifdef AXI_NSPV_M16_AR_QOSARB
  `undef AXI_NSPV_M16_AR_QOSARB
`endif 

`ifdef AXI_NSPV_M1_AW_QOSARB
  `undef AXI_NSPV_M1_AW_QOSARB
`endif 

`ifdef AXI_NSPV_M2_AW_QOSARB
  `undef AXI_NSPV_M2_AW_QOSARB
`endif 

`ifdef AXI_NSPV_M3_AW_QOSARB
  `undef AXI_NSPV_M3_AW_QOSARB
`endif 

`ifdef AXI_NSPV_M4_AW_QOSARB
  `undef AXI_NSPV_M4_AW_QOSARB
`endif 

`ifdef AXI_NSPV_M5_AW_QOSARB
  `undef AXI_NSPV_M5_AW_QOSARB
`endif 

`ifdef AXI_NSPV_M6_AW_QOSARB
  `undef AXI_NSPV_M6_AW_QOSARB
`endif 

`ifdef AXI_NSPV_M7_AW_QOSARB
  `undef AXI_NSPV_M7_AW_QOSARB
`endif 

`ifdef AXI_NSPV_M8_AW_QOSARB
  `undef AXI_NSPV_M8_AW_QOSARB
`endif 

`ifdef AXI_NSPV_M9_AW_QOSARB
  `undef AXI_NSPV_M9_AW_QOSARB
`endif 

`ifdef AXI_NSPV_M10_AW_QOSARB
  `undef AXI_NSPV_M10_AW_QOSARB
`endif 

`ifdef AXI_NSPV_M11_AW_QOSARB
  `undef AXI_NSPV_M11_AW_QOSARB
`endif 

`ifdef AXI_NSPV_M12_AW_QOSARB
  `undef AXI_NSPV_M12_AW_QOSARB
`endif 

`ifdef AXI_NSPV_M13_AW_QOSARB
  `undef AXI_NSPV_M13_AW_QOSARB
`endif 

`ifdef AXI_NSPV_M14_AW_QOSARB
  `undef AXI_NSPV_M14_AW_QOSARB
`endif 

`ifdef AXI_NSPV_M15_AW_QOSARB
  `undef AXI_NSPV_M15_AW_QOSARB
`endif 

`ifdef AXI_NSPV_M16_AW_QOSARB
  `undef AXI_NSPV_M16_AW_QOSARB
`endif 

`ifdef AXI_AR_HAS_QOS_REGULATOR_M1
  `undef AXI_AR_HAS_QOS_REGULATOR_M1
`endif 

`ifdef AXI_AR_QOS_REGULATOR_M1
  `undef AXI_AR_QOS_REGULATOR_M1
`endif 

`ifdef AXI_AR_HAS_QOS_REGULATOR_M2
  `undef AXI_AR_HAS_QOS_REGULATOR_M2
`endif 

`ifdef AXI_AR_QOS_REGULATOR_M2
  `undef AXI_AR_QOS_REGULATOR_M2
`endif 

`ifdef AXI_AR_HAS_QOS_REGULATOR_M3
  `undef AXI_AR_HAS_QOS_REGULATOR_M3
`endif 

`ifdef AXI_AR_QOS_REGULATOR_M3
  `undef AXI_AR_QOS_REGULATOR_M3
`endif 

`ifdef AXI_AR_HAS_QOS_REGULATOR_M4
  `undef AXI_AR_HAS_QOS_REGULATOR_M4
`endif 

`ifdef AXI_AR_QOS_REGULATOR_M4
  `undef AXI_AR_QOS_REGULATOR_M4
`endif 

`ifdef AXI_AR_HAS_QOS_REGULATOR_M5
  `undef AXI_AR_HAS_QOS_REGULATOR_M5
`endif 

`ifdef AXI_AR_QOS_REGULATOR_M5
  `undef AXI_AR_QOS_REGULATOR_M5
`endif 

`ifdef AXI_AR_HAS_QOS_REGULATOR_M6
  `undef AXI_AR_HAS_QOS_REGULATOR_M6
`endif 

`ifdef AXI_AR_QOS_REGULATOR_M6
  `undef AXI_AR_QOS_REGULATOR_M6
`endif 

`ifdef AXI_AR_HAS_QOS_REGULATOR_M7
  `undef AXI_AR_HAS_QOS_REGULATOR_M7
`endif 

`ifdef AXI_AR_QOS_REGULATOR_M7
  `undef AXI_AR_QOS_REGULATOR_M7
`endif 

`ifdef AXI_AR_HAS_QOS_REGULATOR_M8
  `undef AXI_AR_HAS_QOS_REGULATOR_M8
`endif 

`ifdef AXI_AR_QOS_REGULATOR_M8
  `undef AXI_AR_QOS_REGULATOR_M8
`endif 

`ifdef AXI_AR_HAS_QOS_REGULATOR_M9
  `undef AXI_AR_HAS_QOS_REGULATOR_M9
`endif 

`ifdef AXI_AR_QOS_REGULATOR_M9
  `undef AXI_AR_QOS_REGULATOR_M9
`endif 

`ifdef AXI_AR_HAS_QOS_REGULATOR_M10
  `undef AXI_AR_HAS_QOS_REGULATOR_M10
`endif 

`ifdef AXI_AR_QOS_REGULATOR_M10
  `undef AXI_AR_QOS_REGULATOR_M10
`endif 

`ifdef AXI_AR_HAS_QOS_REGULATOR_M11
  `undef AXI_AR_HAS_QOS_REGULATOR_M11
`endif 

`ifdef AXI_AR_QOS_REGULATOR_M11
  `undef AXI_AR_QOS_REGULATOR_M11
`endif 

`ifdef AXI_AR_HAS_QOS_REGULATOR_M12
  `undef AXI_AR_HAS_QOS_REGULATOR_M12
`endif 

`ifdef AXI_AR_QOS_REGULATOR_M12
  `undef AXI_AR_QOS_REGULATOR_M12
`endif 

`ifdef AXI_AR_HAS_QOS_REGULATOR_M13
  `undef AXI_AR_HAS_QOS_REGULATOR_M13
`endif 

`ifdef AXI_AR_QOS_REGULATOR_M13
  `undef AXI_AR_QOS_REGULATOR_M13
`endif 

`ifdef AXI_AR_HAS_QOS_REGULATOR_M14
  `undef AXI_AR_HAS_QOS_REGULATOR_M14
`endif 

`ifdef AXI_AR_QOS_REGULATOR_M14
  `undef AXI_AR_QOS_REGULATOR_M14
`endif 

`ifdef AXI_AR_HAS_QOS_REGULATOR_M15
  `undef AXI_AR_HAS_QOS_REGULATOR_M15
`endif 

`ifdef AXI_AR_QOS_REGULATOR_M15
  `undef AXI_AR_QOS_REGULATOR_M15
`endif 

`ifdef AXI_AR_HAS_QOS_REGULATOR_M16
  `undef AXI_AR_HAS_QOS_REGULATOR_M16
`endif 

`ifdef AXI_AR_QOS_REGULATOR_M16
  `undef AXI_AR_QOS_REGULATOR_M16
`endif 

`ifdef AXI_AW_HAS_QOS_REGULATOR_M1
  `undef AXI_AW_HAS_QOS_REGULATOR_M1
`endif 

`ifdef AXI_AW_QOS_REGULATOR_M1
  `undef AXI_AW_QOS_REGULATOR_M1
`endif 

`ifdef AXI_AW_HAS_QOS_REGULATOR_M2
  `undef AXI_AW_HAS_QOS_REGULATOR_M2
`endif 

`ifdef AXI_AW_QOS_REGULATOR_M2
  `undef AXI_AW_QOS_REGULATOR_M2
`endif 

`ifdef AXI_AW_HAS_QOS_REGULATOR_M3
  `undef AXI_AW_HAS_QOS_REGULATOR_M3
`endif 

`ifdef AXI_AW_QOS_REGULATOR_M3
  `undef AXI_AW_QOS_REGULATOR_M3
`endif 

`ifdef AXI_AW_HAS_QOS_REGULATOR_M4
  `undef AXI_AW_HAS_QOS_REGULATOR_M4
`endif 

`ifdef AXI_AW_QOS_REGULATOR_M4
  `undef AXI_AW_QOS_REGULATOR_M4
`endif 

`ifdef AXI_AW_HAS_QOS_REGULATOR_M5
  `undef AXI_AW_HAS_QOS_REGULATOR_M5
`endif 

`ifdef AXI_AW_QOS_REGULATOR_M5
  `undef AXI_AW_QOS_REGULATOR_M5
`endif 

`ifdef AXI_AW_HAS_QOS_REGULATOR_M6
  `undef AXI_AW_HAS_QOS_REGULATOR_M6
`endif 

`ifdef AXI_AW_QOS_REGULATOR_M6
  `undef AXI_AW_QOS_REGULATOR_M6
`endif 

`ifdef AXI_AW_HAS_QOS_REGULATOR_M7
  `undef AXI_AW_HAS_QOS_REGULATOR_M7
`endif 

`ifdef AXI_AW_QOS_REGULATOR_M7
  `undef AXI_AW_QOS_REGULATOR_M7
`endif 

`ifdef AXI_AW_HAS_QOS_REGULATOR_M8
  `undef AXI_AW_HAS_QOS_REGULATOR_M8
`endif 

`ifdef AXI_AW_QOS_REGULATOR_M8
  `undef AXI_AW_QOS_REGULATOR_M8
`endif 

`ifdef AXI_AW_HAS_QOS_REGULATOR_M9
  `undef AXI_AW_HAS_QOS_REGULATOR_M9
`endif 

`ifdef AXI_AW_QOS_REGULATOR_M9
  `undef AXI_AW_QOS_REGULATOR_M9
`endif 

`ifdef AXI_AW_HAS_QOS_REGULATOR_M10
  `undef AXI_AW_HAS_QOS_REGULATOR_M10
`endif 

`ifdef AXI_AW_QOS_REGULATOR_M10
  `undef AXI_AW_QOS_REGULATOR_M10
`endif 

`ifdef AXI_AW_HAS_QOS_REGULATOR_M11
  `undef AXI_AW_HAS_QOS_REGULATOR_M11
`endif 

`ifdef AXI_AW_QOS_REGULATOR_M11
  `undef AXI_AW_QOS_REGULATOR_M11
`endif 

`ifdef AXI_AW_HAS_QOS_REGULATOR_M12
  `undef AXI_AW_HAS_QOS_REGULATOR_M12
`endif 

`ifdef AXI_AW_QOS_REGULATOR_M12
  `undef AXI_AW_QOS_REGULATOR_M12
`endif 

`ifdef AXI_AW_HAS_QOS_REGULATOR_M13
  `undef AXI_AW_HAS_QOS_REGULATOR_M13
`endif 

`ifdef AXI_AW_QOS_REGULATOR_M13
  `undef AXI_AW_QOS_REGULATOR_M13
`endif 

`ifdef AXI_AW_HAS_QOS_REGULATOR_M14
  `undef AXI_AW_HAS_QOS_REGULATOR_M14
`endif 

`ifdef AXI_AW_QOS_REGULATOR_M14
  `undef AXI_AW_QOS_REGULATOR_M14
`endif 

`ifdef AXI_AW_HAS_QOS_REGULATOR_M15
  `undef AXI_AW_HAS_QOS_REGULATOR_M15
`endif 

`ifdef AXI_AW_QOS_REGULATOR_M15
  `undef AXI_AW_QOS_REGULATOR_M15
`endif 

`ifdef AXI_AW_HAS_QOS_REGULATOR_M16
  `undef AXI_AW_HAS_QOS_REGULATOR_M16
`endif 

`ifdef AXI_AW_QOS_REGULATOR_M16
  `undef AXI_AW_QOS_REGULATOR_M16
`endif 

`ifdef AXI_HAS_ARQOS_EXT_M1
  `undef AXI_HAS_ARQOS_EXT_M1
`endif 

`ifdef AXI_ARQOS_EXT_M1
  `undef AXI_ARQOS_EXT_M1
`endif 

`ifdef AXI_ARQOS_INT_M1
  `undef AXI_ARQOS_INT_M1
`endif 

`ifdef AXI_HAS_ARQOS_EXT_M2
  `undef AXI_HAS_ARQOS_EXT_M2
`endif 

`ifdef AXI_ARQOS_EXT_M2
  `undef AXI_ARQOS_EXT_M2
`endif 

`ifdef AXI_ARQOS_INT_M2
  `undef AXI_ARQOS_INT_M2
`endif 

`ifdef AXI_HAS_ARQOS_EXT_M3
  `undef AXI_HAS_ARQOS_EXT_M3
`endif 

`ifdef AXI_ARQOS_EXT_M3
  `undef AXI_ARQOS_EXT_M3
`endif 

`ifdef AXI_ARQOS_INT_M3
  `undef AXI_ARQOS_INT_M3
`endif 

`ifdef AXI_HAS_ARQOS_EXT_M4
  `undef AXI_HAS_ARQOS_EXT_M4
`endif 

`ifdef AXI_ARQOS_EXT_M4
  `undef AXI_ARQOS_EXT_M4
`endif 

`ifdef AXI_ARQOS_INT_M4
  `undef AXI_ARQOS_INT_M4
`endif 

`ifdef AXI_HAS_ARQOS_EXT_M5
  `undef AXI_HAS_ARQOS_EXT_M5
`endif 

`ifdef AXI_ARQOS_EXT_M5
  `undef AXI_ARQOS_EXT_M5
`endif 

`ifdef AXI_ARQOS_INT_M5
  `undef AXI_ARQOS_INT_M5
`endif 

`ifdef AXI_HAS_ARQOS_EXT_M6
  `undef AXI_HAS_ARQOS_EXT_M6
`endif 

`ifdef AXI_ARQOS_EXT_M6
  `undef AXI_ARQOS_EXT_M6
`endif 

`ifdef AXI_ARQOS_INT_M6
  `undef AXI_ARQOS_INT_M6
`endif 

`ifdef AXI_HAS_ARQOS_EXT_M7
  `undef AXI_HAS_ARQOS_EXT_M7
`endif 

`ifdef AXI_ARQOS_EXT_M7
  `undef AXI_ARQOS_EXT_M7
`endif 

`ifdef AXI_ARQOS_INT_M7
  `undef AXI_ARQOS_INT_M7
`endif 

`ifdef AXI_HAS_ARQOS_EXT_M8
  `undef AXI_HAS_ARQOS_EXT_M8
`endif 

`ifdef AXI_ARQOS_EXT_M8
  `undef AXI_ARQOS_EXT_M8
`endif 

`ifdef AXI_ARQOS_INT_M8
  `undef AXI_ARQOS_INT_M8
`endif 

`ifdef AXI_HAS_ARQOS_EXT_M9
  `undef AXI_HAS_ARQOS_EXT_M9
`endif 

`ifdef AXI_ARQOS_EXT_M9
  `undef AXI_ARQOS_EXT_M9
`endif 

`ifdef AXI_ARQOS_INT_M9
  `undef AXI_ARQOS_INT_M9
`endif 

`ifdef AXI_HAS_ARQOS_EXT_M10
  `undef AXI_HAS_ARQOS_EXT_M10
`endif 

`ifdef AXI_ARQOS_EXT_M10
  `undef AXI_ARQOS_EXT_M10
`endif 

`ifdef AXI_ARQOS_INT_M10
  `undef AXI_ARQOS_INT_M10
`endif 

`ifdef AXI_HAS_ARQOS_EXT_M11
  `undef AXI_HAS_ARQOS_EXT_M11
`endif 

`ifdef AXI_ARQOS_EXT_M11
  `undef AXI_ARQOS_EXT_M11
`endif 

`ifdef AXI_ARQOS_INT_M11
  `undef AXI_ARQOS_INT_M11
`endif 

`ifdef AXI_HAS_ARQOS_EXT_M12
  `undef AXI_HAS_ARQOS_EXT_M12
`endif 

`ifdef AXI_ARQOS_EXT_M12
  `undef AXI_ARQOS_EXT_M12
`endif 

`ifdef AXI_ARQOS_INT_M12
  `undef AXI_ARQOS_INT_M12
`endif 

`ifdef AXI_HAS_ARQOS_EXT_M13
  `undef AXI_HAS_ARQOS_EXT_M13
`endif 

`ifdef AXI_ARQOS_EXT_M13
  `undef AXI_ARQOS_EXT_M13
`endif 

`ifdef AXI_ARQOS_INT_M13
  `undef AXI_ARQOS_INT_M13
`endif 

`ifdef AXI_HAS_ARQOS_EXT_M14
  `undef AXI_HAS_ARQOS_EXT_M14
`endif 

`ifdef AXI_ARQOS_EXT_M14
  `undef AXI_ARQOS_EXT_M14
`endif 

`ifdef AXI_ARQOS_INT_M14
  `undef AXI_ARQOS_INT_M14
`endif 

`ifdef AXI_HAS_ARQOS_EXT_M15
  `undef AXI_HAS_ARQOS_EXT_M15
`endif 

`ifdef AXI_ARQOS_EXT_M15
  `undef AXI_ARQOS_EXT_M15
`endif 

`ifdef AXI_ARQOS_INT_M15
  `undef AXI_ARQOS_INT_M15
`endif 

`ifdef AXI_HAS_ARQOS_EXT_M16
  `undef AXI_HAS_ARQOS_EXT_M16
`endif 

`ifdef AXI_ARQOS_EXT_M16
  `undef AXI_ARQOS_EXT_M16
`endif 

`ifdef AXI_ARQOS_INT_M16
  `undef AXI_ARQOS_INT_M16
`endif 

`ifdef AXI_HAS_AWQOS_EXT_M1
  `undef AXI_HAS_AWQOS_EXT_M1
`endif 

`ifdef AXI_AWQOS_EXT_M1
  `undef AXI_AWQOS_EXT_M1
`endif 

`ifdef AXI_AWQOS_INT_M1
  `undef AXI_AWQOS_INT_M1
`endif 

`ifdef AXI_HAS_AWQOS_EXT_M2
  `undef AXI_HAS_AWQOS_EXT_M2
`endif 

`ifdef AXI_AWQOS_EXT_M2
  `undef AXI_AWQOS_EXT_M2
`endif 

`ifdef AXI_AWQOS_INT_M2
  `undef AXI_AWQOS_INT_M2
`endif 

`ifdef AXI_HAS_AWQOS_EXT_M3
  `undef AXI_HAS_AWQOS_EXT_M3
`endif 

`ifdef AXI_AWQOS_EXT_M3
  `undef AXI_AWQOS_EXT_M3
`endif 

`ifdef AXI_AWQOS_INT_M3
  `undef AXI_AWQOS_INT_M3
`endif 

`ifdef AXI_HAS_AWQOS_EXT_M4
  `undef AXI_HAS_AWQOS_EXT_M4
`endif 

`ifdef AXI_AWQOS_EXT_M4
  `undef AXI_AWQOS_EXT_M4
`endif 

`ifdef AXI_AWQOS_INT_M4
  `undef AXI_AWQOS_INT_M4
`endif 

`ifdef AXI_HAS_AWQOS_EXT_M5
  `undef AXI_HAS_AWQOS_EXT_M5
`endif 

`ifdef AXI_AWQOS_EXT_M5
  `undef AXI_AWQOS_EXT_M5
`endif 

`ifdef AXI_AWQOS_INT_M5
  `undef AXI_AWQOS_INT_M5
`endif 

`ifdef AXI_HAS_AWQOS_EXT_M6
  `undef AXI_HAS_AWQOS_EXT_M6
`endif 

`ifdef AXI_AWQOS_EXT_M6
  `undef AXI_AWQOS_EXT_M6
`endif 

`ifdef AXI_AWQOS_INT_M6
  `undef AXI_AWQOS_INT_M6
`endif 

`ifdef AXI_HAS_AWQOS_EXT_M7
  `undef AXI_HAS_AWQOS_EXT_M7
`endif 

`ifdef AXI_AWQOS_EXT_M7
  `undef AXI_AWQOS_EXT_M7
`endif 

`ifdef AXI_AWQOS_INT_M7
  `undef AXI_AWQOS_INT_M7
`endif 

`ifdef AXI_HAS_AWQOS_EXT_M8
  `undef AXI_HAS_AWQOS_EXT_M8
`endif 

`ifdef AXI_AWQOS_EXT_M8
  `undef AXI_AWQOS_EXT_M8
`endif 

`ifdef AXI_AWQOS_INT_M8
  `undef AXI_AWQOS_INT_M8
`endif 

`ifdef AXI_HAS_AWQOS_EXT_M9
  `undef AXI_HAS_AWQOS_EXT_M9
`endif 

`ifdef AXI_AWQOS_EXT_M9
  `undef AXI_AWQOS_EXT_M9
`endif 

`ifdef AXI_AWQOS_INT_M9
  `undef AXI_AWQOS_INT_M9
`endif 

`ifdef AXI_HAS_AWQOS_EXT_M10
  `undef AXI_HAS_AWQOS_EXT_M10
`endif 

`ifdef AXI_AWQOS_EXT_M10
  `undef AXI_AWQOS_EXT_M10
`endif 

`ifdef AXI_AWQOS_INT_M10
  `undef AXI_AWQOS_INT_M10
`endif 

`ifdef AXI_HAS_AWQOS_EXT_M11
  `undef AXI_HAS_AWQOS_EXT_M11
`endif 

`ifdef AXI_AWQOS_EXT_M11
  `undef AXI_AWQOS_EXT_M11
`endif 

`ifdef AXI_AWQOS_INT_M11
  `undef AXI_AWQOS_INT_M11
`endif 

`ifdef AXI_HAS_AWQOS_EXT_M12
  `undef AXI_HAS_AWQOS_EXT_M12
`endif 

`ifdef AXI_AWQOS_EXT_M12
  `undef AXI_AWQOS_EXT_M12
`endif 

`ifdef AXI_AWQOS_INT_M12
  `undef AXI_AWQOS_INT_M12
`endif 

`ifdef AXI_HAS_AWQOS_EXT_M13
  `undef AXI_HAS_AWQOS_EXT_M13
`endif 

`ifdef AXI_AWQOS_EXT_M13
  `undef AXI_AWQOS_EXT_M13
`endif 

`ifdef AXI_AWQOS_INT_M13
  `undef AXI_AWQOS_INT_M13
`endif 

`ifdef AXI_HAS_AWQOS_EXT_M14
  `undef AXI_HAS_AWQOS_EXT_M14
`endif 

`ifdef AXI_AWQOS_EXT_M14
  `undef AXI_AWQOS_EXT_M14
`endif 

`ifdef AXI_AWQOS_INT_M14
  `undef AXI_AWQOS_INT_M14
`endif 

`ifdef AXI_HAS_AWQOS_EXT_M15
  `undef AXI_HAS_AWQOS_EXT_M15
`endif 

`ifdef AXI_AWQOS_EXT_M15
  `undef AXI_AWQOS_EXT_M15
`endif 

`ifdef AXI_AWQOS_INT_M15
  `undef AXI_AWQOS_INT_M15
`endif 

`ifdef AXI_HAS_AWQOS_EXT_M16
  `undef AXI_HAS_AWQOS_EXT_M16
`endif 

`ifdef AXI_AWQOS_EXT_M16
  `undef AXI_AWQOS_EXT_M16
`endif 

`ifdef AXI_AWQOS_INT_M16
  `undef AXI_AWQOS_INT_M16
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AR_S0
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AR_S0
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AR_S1
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AR_S1
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AR_S2
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AR_S2
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AR_S3
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AR_S3
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AR_S4
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AR_S4
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AR_S5
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AR_S5
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AR_S6
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AR_S6
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AR_S7
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AR_S7
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AR_S8
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AR_S8
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AR_S9
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AR_S9
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AR_S10
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AR_S10
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AR_S11
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AR_S11
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AR_S12
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AR_S12
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AR_S13
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AR_S13
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AR_S14
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AR_S14
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AR_S15
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AR_S15
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AR_S16
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AR_S16
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AW_S0
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AW_S0
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AW_S1
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AW_S1
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AW_S2
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AW_S2
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AW_S3
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AW_S3
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AW_S4
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AW_S4
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AW_S5
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AW_S5
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AW_S6
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AW_S6
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AW_S7
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AW_S7
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AW_S8
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AW_S8
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AW_S9
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AW_S9
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AW_S10
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AW_S10
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AW_S11
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AW_S11
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AW_S12
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AW_S12
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AW_S13
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AW_S13
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AW_S14
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AW_S14
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AW_S15
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AW_S15
`endif 

`ifdef AXI_HAS_QOS_ARB_TYPE_ON_AW_S16
  `undef AXI_HAS_QOS_ARB_TYPE_ON_AW_S16
`endif 

`ifdef SNPS_RCE_INTERNAL_ON
  `undef SNPS_RCE_INTERNAL_ON
`endif 

`ifdef AXI_DW_GT_64
  `undef AXI_DW_GT_64
`endif 

`ifdef AXI_HAS_APB
  `undef AXI_HAS_APB
`endif 

`ifdef AXI_HAS_APB3
  `undef AXI_HAS_APB3
`endif 

`ifdef AXI_APB3
  `undef AXI_APB3
`endif 

`ifdef APB_DATA_WIDTH
  `undef APB_DATA_WIDTH
`endif 

`ifdef AXI_IC_REG_BASE_ADDR
  `undef AXI_IC_REG_BASE_ADDR
`endif 

`ifdef AXI_NUM_SYNC_FF
  `undef AXI_NUM_SYNC_FF
`endif 

`ifdef DW_AXI_VERSION_ID
  `undef DW_AXI_VERSION_ID
`endif 

`ifdef AXI_VERIF_EN
  `undef AXI_VERIF_EN
`endif 

`ifdef AXI_4
  `undef AXI_4
`endif 

`ifdef AXI_ACELITE
  `undef AXI_ACELITE
`endif 

`ifdef AXI_HAS_REGIONS_S1
  `undef AXI_HAS_REGIONS_S1
`endif 

`ifdef AXI_REGIONS_S1
  `undef AXI_REGIONS_S1
`endif 

`ifdef AXI_HAS_REGIONS_S2
  `undef AXI_HAS_REGIONS_S2
`endif 

`ifdef AXI_REGIONS_S2
  `undef AXI_REGIONS_S2
`endif 

`ifdef AXI_HAS_REGIONS_S3
  `undef AXI_HAS_REGIONS_S3
`endif 

`ifdef AXI_REGIONS_S3
  `undef AXI_REGIONS_S3
`endif 

`ifdef AXI_HAS_REGIONS_S4
  `undef AXI_HAS_REGIONS_S4
`endif 

`ifdef AXI_REGIONS_S4
  `undef AXI_REGIONS_S4
`endif 

`ifdef AXI_HAS_REGIONS_S5
  `undef AXI_HAS_REGIONS_S5
`endif 

`ifdef AXI_REGIONS_S5
  `undef AXI_REGIONS_S5
`endif 

`ifdef AXI_HAS_REGIONS_S6
  `undef AXI_HAS_REGIONS_S6
`endif 

`ifdef AXI_REGIONS_S6
  `undef AXI_REGIONS_S6
`endif 

`ifdef AXI_HAS_REGIONS_S7
  `undef AXI_HAS_REGIONS_S7
`endif 

`ifdef AXI_REGIONS_S7
  `undef AXI_REGIONS_S7
`endif 

`ifdef AXI_HAS_REGIONS_S8
  `undef AXI_HAS_REGIONS_S8
`endif 

`ifdef AXI_REGIONS_S8
  `undef AXI_REGIONS_S8
`endif 

`ifdef AXI_HAS_REGIONS_S9
  `undef AXI_HAS_REGIONS_S9
`endif 

`ifdef AXI_REGIONS_S9
  `undef AXI_REGIONS_S9
`endif 

`ifdef AXI_HAS_REGIONS_S10
  `undef AXI_HAS_REGIONS_S10
`endif 

`ifdef AXI_REGIONS_S10
  `undef AXI_REGIONS_S10
`endif 

`ifdef AXI_HAS_REGIONS_S11
  `undef AXI_HAS_REGIONS_S11
`endif 

`ifdef AXI_REGIONS_S11
  `undef AXI_REGIONS_S11
`endif 

`ifdef AXI_HAS_REGIONS_S12
  `undef AXI_HAS_REGIONS_S12
`endif 

`ifdef AXI_REGIONS_S12
  `undef AXI_REGIONS_S12
`endif 

`ifdef AXI_HAS_REGIONS_S13
  `undef AXI_HAS_REGIONS_S13
`endif 

`ifdef AXI_REGIONS_S13
  `undef AXI_REGIONS_S13
`endif 

`ifdef AXI_HAS_REGIONS_S14
  `undef AXI_HAS_REGIONS_S14
`endif 

`ifdef AXI_REGIONS_S14
  `undef AXI_REGIONS_S14
`endif 

`ifdef AXI_HAS_REGIONS_S15
  `undef AXI_HAS_REGIONS_S15
`endif 

`ifdef AXI_REGIONS_S15
  `undef AXI_REGIONS_S15
`endif 

`ifdef AXI_HAS_REGIONS_S16
  `undef AXI_HAS_REGIONS_S16
`endif 

`ifdef AXI_REGIONS_S16
  `undef AXI_REGIONS_S16
`endif 

`ifdef AXI_HAS_REGIONS
  `undef AXI_HAS_REGIONS
`endif 

`ifdef AXI_REGIONS
  `undef AXI_REGIONS
`endif 

`ifdef AXI_LEGACY_LP_MODE
  `undef AXI_LEGACY_LP_MODE
`endif 

`ifdef AXI_BCM_TST_MODE
  `undef AXI_BCM_TST_MODE
`endif 

`ifdef AXI_BCM_CDC_INIT
  `undef AXI_BCM_CDC_INIT
`endif 

`ifdef DWC_NO_TST_MODE
  `undef DWC_NO_TST_MODE
`endif 

`ifdef DWC_NO_CDC_INIT
  `undef DWC_NO_CDC_INIT
`endif 

`ifdef __GUARD__DW_AXI_CONSTANTS__VH__
  `undef __GUARD__DW_AXI_CONSTANTS__VH__
`endif 

`ifdef AXI_BSW
  `undef AXI_BSW
`endif 

`ifdef AXI_BTW
  `undef AXI_BTW
`endif 

`ifdef AXI_LTW
  `undef AXI_LTW
`endif 

`ifdef AXI_CTW
  `undef AXI_CTW
`endif 

`ifdef AXI_PTW
  `undef AXI_PTW
`endif 

`ifdef AXI_BRW
  `undef AXI_BRW
`endif 

`ifdef AXI_RRW
  `undef AXI_RRW
`endif 

`ifdef AXI_SW
  `undef AXI_SW
`endif 

`ifdef AXI_MAX_NUM_MST_SLVS
  `undef AXI_MAX_NUM_MST_SLVS
`endif 

`ifdef AXI_MAX_NUM_USR_MSTS
  `undef AXI_MAX_NUM_USR_MSTS
`endif 

`ifdef AXI_MAX_NUM_USR_SLVS
  `undef AXI_MAX_NUM_USR_SLVS
`endif 

`ifdef AXI_LT_NORM
  `undef AXI_LT_NORM
`endif 

`ifdef AXI_LT_EX
  `undef AXI_LT_EX
`endif 

`ifdef AXI_LT_LOCK
  `undef AXI_LT_LOCK
`endif 

`ifdef AXI_PT_PRVLGD
  `undef AXI_PT_PRVLGD
`endif 

`ifdef AXI_PT_NORM
  `undef AXI_PT_NORM
`endif 

`ifdef AXI_PT_SECURE
  `undef AXI_PT_SECURE
`endif 

`ifdef AXI_PT_NSECURE
  `undef AXI_PT_NSECURE
`endif 

`ifdef AXI_PT_INSTRUCT
  `undef AXI_PT_INSTRUCT
`endif 

`ifdef AXI_PT_DATA
  `undef AXI_PT_DATA
`endif 

`ifdef AXI_PT_PRVLGD_BIT
  `undef AXI_PT_PRVLGD_BIT
`endif 

`ifdef AXI_PT_INSTRUCT_BIT
  `undef AXI_PT_INSTRUCT_BIT
`endif 

`ifdef AXI_RESP_OKAY
  `undef AXI_RESP_OKAY
`endif 

`ifdef AXI_RESP_EXOKAY
  `undef AXI_RESP_EXOKAY
`endif 

`ifdef AXI_RESP_SLVERR
  `undef AXI_RESP_SLVERR
`endif 

`ifdef AXI_RESP_DECERR
  `undef AXI_RESP_DECERR
`endif 

`ifdef AXI_TMO_COMB
  `undef AXI_TMO_COMB
`endif 

`ifdef AXI_TMO_FRWD
  `undef AXI_TMO_FRWD
`endif 

`ifdef AXI_TMO_FULL
  `undef AXI_TMO_FULL
`endif 

`ifdef AXI_NOREQ_LOCKING
  `undef AXI_NOREQ_LOCKING
`endif 

`ifdef AXI_REQ_LOCKING
  `undef AXI_REQ_LOCKING
`endif 

`ifdef AXI_ARB_TYPE_DP
  `undef AXI_ARB_TYPE_DP
`endif 

`ifdef AXI_ARB_TYPE_FCFS
  `undef AXI_ARB_TYPE_FCFS
`endif 

`ifdef AXI_ARB_TYPE_2T
  `undef AXI_ARB_TYPE_2T
`endif 

`ifdef AXI_ARB_TYPE_USER
  `undef AXI_ARB_TYPE_USER
`endif 

`ifdef AXI_ARB_TYPE_QOS
  `undef AXI_ARB_TYPE_QOS
`endif 

`ifdef AXI_W_CH
  `undef AXI_W_CH
`endif 

`ifdef AXI_NOT_W_CH
  `undef AXI_NOT_W_CH
`endif 

`ifdef AXI_AW_CH
  `undef AXI_AW_CH
`endif 

`ifdef AXI_NOT_AW_CH
  `undef AXI_NOT_AW_CH
`endif 

`ifdef AXI_R_CH
  `undef AXI_R_CH
`endif 

`ifdef AXI_NOT_R_CH
  `undef AXI_NOT_R_CH
`endif 

`ifdef AXI_ADDR_CH
  `undef AXI_ADDR_CH
`endif 

`ifdef AXI_NOT_ADDR_CH
  `undef AXI_NOT_ADDR_CH
`endif 

`ifdef USE_INT_GI
  `undef USE_INT_GI
`endif 

`ifdef USE_EXT_GI
  `undef USE_EXT_GI
`endif 

`ifdef AXI_SHARED
  `undef AXI_SHARED
`endif 

`ifdef AXI_NOT_SHARED
  `undef AXI_NOT_SHARED
`endif 

`ifdef AXI_HOLD_VLD_OTHER_S_W
  `undef AXI_HOLD_VLD_OTHER_S_W
`endif 

`ifdef AXI_HOLD_VLD_OTHER_M_W
  `undef AXI_HOLD_VLD_OTHER_M_W
`endif 

`ifdef AXI_ARPYLD_PROT_RHS
  `undef AXI_ARPYLD_PROT_RHS
`endif 

`ifdef AXI_ARPYLD_PROT_LHS
  `undef AXI_ARPYLD_PROT_LHS
`endif 

`ifdef AXI_ARPYLD_PROT
  `undef AXI_ARPYLD_PROT
`endif 

`ifdef AXI_ARPYLD_CACHE_RHS
  `undef AXI_ARPYLD_CACHE_RHS
`endif 

`ifdef AXI_ARPYLD_CACHE_LHS
  `undef AXI_ARPYLD_CACHE_LHS
`endif 

`ifdef AXI_ARPYLD_CACHE
  `undef AXI_ARPYLD_CACHE
`endif 

`ifdef AXI_ARPYLD_LOCK_RHS
  `undef AXI_ARPYLD_LOCK_RHS
`endif 

`ifdef AXI_ARPYLD_LOCK_LHS
  `undef AXI_ARPYLD_LOCK_LHS
`endif 

`ifdef AXI_ARPYLD_LOCK
  `undef AXI_ARPYLD_LOCK
`endif 

`ifdef AXI_ARPYLD_BURST_RHS
  `undef AXI_ARPYLD_BURST_RHS
`endif 

`ifdef AXI_ARPYLD_BURST_LHS
  `undef AXI_ARPYLD_BURST_LHS
`endif 

`ifdef AXI_ARPYLD_BURST
  `undef AXI_ARPYLD_BURST
`endif 

`ifdef AXI_ARPYLD_SIZE_RHS
  `undef AXI_ARPYLD_SIZE_RHS
`endif 

`ifdef AXI_ARPYLD_SIZE_LHS
  `undef AXI_ARPYLD_SIZE_LHS
`endif 

`ifdef AXI_ARPYLD_SIZE
  `undef AXI_ARPYLD_SIZE
`endif 

`ifdef AXI_ARPYLD_LEN_RHS
  `undef AXI_ARPYLD_LEN_RHS
`endif 

`ifdef AXI_ARPYLD_LEN_LHS
  `undef AXI_ARPYLD_LEN_LHS
`endif 

`ifdef AXI_ARPYLD_LEN
  `undef AXI_ARPYLD_LEN
`endif 

`ifdef AXI_ARPYLD_ADDR_RHS
  `undef AXI_ARPYLD_ADDR_RHS
`endif 

`ifdef AXI_ARPYLD_ADDR_LHS
  `undef AXI_ARPYLD_ADDR_LHS
`endif 

`ifdef AXI_ARPYLD_ADDR
  `undef AXI_ARPYLD_ADDR
`endif 

`ifdef AXI_ARPYLD_ID_RHS_M
  `undef AXI_ARPYLD_ID_RHS_M
`endif 

`ifdef AXI_ARPYLD_ID_LHS_M
  `undef AXI_ARPYLD_ID_LHS_M
`endif 

`ifdef AXI_ARPYLD_ID_M
  `undef AXI_ARPYLD_ID_M
`endif 

`ifdef AXI_ARPYLD_ID_RHS_S
  `undef AXI_ARPYLD_ID_RHS_S
`endif 

`ifdef AXI_ARPYLD_ID_LHS_S
  `undef AXI_ARPYLD_ID_LHS_S
`endif 

`ifdef AXI_ARPYLD_ID_S
  `undef AXI_ARPYLD_ID_S
`endif 

`ifdef AXI_RPYLD_LAST_LHS
  `undef AXI_RPYLD_LAST_LHS
`endif 

`ifdef AXI_RPYLD_LAST
  `undef AXI_RPYLD_LAST
`endif 

`ifdef AXI_RPYLD_RESP_RHS
  `undef AXI_RPYLD_RESP_RHS
`endif 

`ifdef AXI_RPYLD_RESP_LHS
  `undef AXI_RPYLD_RESP_LHS
`endif 

`ifdef AXI_RPYLD_RESP
  `undef AXI_RPYLD_RESP
`endif 

`ifdef AXI_RPYLD_DATA_RHS
  `undef AXI_RPYLD_DATA_RHS
`endif 

`ifdef AXI_RPYLD_DATA_LHS
  `undef AXI_RPYLD_DATA_LHS
`endif 

`ifdef AXI_RPYLD_DATA
  `undef AXI_RPYLD_DATA
`endif 

`ifdef AXI_RPYLD_ID_RHS_M
  `undef AXI_RPYLD_ID_RHS_M
`endif 

`ifdef AXI_RPYLD_ID_LHS_M
  `undef AXI_RPYLD_ID_LHS_M
`endif 

`ifdef AXI_RPYLD_ID_M
  `undef AXI_RPYLD_ID_M
`endif 

`ifdef AXI_RPYLD_ID_RHS_S
  `undef AXI_RPYLD_ID_RHS_S
`endif 

`ifdef AXI_RPYLD_ID_LHS_S
  `undef AXI_RPYLD_ID_LHS_S
`endif 

`ifdef AXI_RPYLD_ID_S
  `undef AXI_RPYLD_ID_S
`endif 

`ifdef AXI_AWPYLD_PROT_RHS
  `undef AXI_AWPYLD_PROT_RHS
`endif 

`ifdef AXI_AWPYLD_PROT_LHS
  `undef AXI_AWPYLD_PROT_LHS
`endif 

`ifdef AXI_AWPYLD_PROT
  `undef AXI_AWPYLD_PROT
`endif 

`ifdef AXI_AWPYLD_CACHE_RHS
  `undef AXI_AWPYLD_CACHE_RHS
`endif 

`ifdef AXI_AWPYLD_CACHE_LHS
  `undef AXI_AWPYLD_CACHE_LHS
`endif 

`ifdef AXI_AWPYLD_CACHE
  `undef AXI_AWPYLD_CACHE
`endif 

`ifdef AXI_AWPYLD_LOCK_RHS
  `undef AXI_AWPYLD_LOCK_RHS
`endif 

`ifdef AXI_AWPYLD_LOCK_LHS
  `undef AXI_AWPYLD_LOCK_LHS
`endif 

`ifdef AXI_AWPYLD_LOCK
  `undef AXI_AWPYLD_LOCK
`endif 

`ifdef AXI_AWPYLD_BURST_RHS
  `undef AXI_AWPYLD_BURST_RHS
`endif 

`ifdef AXI_AWPYLD_BURST_LHS
  `undef AXI_AWPYLD_BURST_LHS
`endif 

`ifdef AXI_AWPYLD_BURST
  `undef AXI_AWPYLD_BURST
`endif 

`ifdef AXI_AWPYLD_SIZE_RHS
  `undef AXI_AWPYLD_SIZE_RHS
`endif 

`ifdef AXI_AWPYLD_SIZE_LHS
  `undef AXI_AWPYLD_SIZE_LHS
`endif 

`ifdef AXI_AWPYLD_SIZE
  `undef AXI_AWPYLD_SIZE
`endif 

`ifdef AXI_AWPYLD_LEN_RHS
  `undef AXI_AWPYLD_LEN_RHS
`endif 

`ifdef AXI_AWPYLD_LEN_LHS
  `undef AXI_AWPYLD_LEN_LHS
`endif 

`ifdef AXI_AWPYLD_LEN
  `undef AXI_AWPYLD_LEN
`endif 

`ifdef AXI_AWPYLD_ADDR_RHS
  `undef AXI_AWPYLD_ADDR_RHS
`endif 

`ifdef AXI_AWPYLD_ADDR_LHS
  `undef AXI_AWPYLD_ADDR_LHS
`endif 

`ifdef AXI_AWPYLD_ADDR
  `undef AXI_AWPYLD_ADDR
`endif 

`ifdef AXI_AWPYLD_ID_RHS_M
  `undef AXI_AWPYLD_ID_RHS_M
`endif 

`ifdef AXI_AWPYLD_ID_LHS_M
  `undef AXI_AWPYLD_ID_LHS_M
`endif 

`ifdef AXI_AWPYLD_ID_M
  `undef AXI_AWPYLD_ID_M
`endif 

`ifdef AXI_AWPYLD_ID_RHS_S
  `undef AXI_AWPYLD_ID_RHS_S
`endif 

`ifdef AXI_AWPYLD_ID_LHS_S
  `undef AXI_AWPYLD_ID_LHS_S
`endif 

`ifdef AXI_AWPYLD_ID_S
  `undef AXI_AWPYLD_ID_S
`endif 

`ifdef AXI_WPYLD_LAST_LHS
  `undef AXI_WPYLD_LAST_LHS
`endif 

`ifdef AXI_WPYLD_LAST
  `undef AXI_WPYLD_LAST
`endif 

`ifdef AXI_WPYLD_STRB_RHS
  `undef AXI_WPYLD_STRB_RHS
`endif 

`ifdef AXI_WPYLD_STRB_LHS
  `undef AXI_WPYLD_STRB_LHS
`endif 

`ifdef AXI_WPYLD_STRB
  `undef AXI_WPYLD_STRB
`endif 

`ifdef AXI_WPYLD_DATA_RHS
  `undef AXI_WPYLD_DATA_RHS
`endif 

`ifdef AXI_WPYLD_DATA_LHS
  `undef AXI_WPYLD_DATA_LHS
`endif 

`ifdef AXI_WPYLD_DATA
  `undef AXI_WPYLD_DATA
`endif 

`ifdef AXI_WPYLD_ID_RHS_M
  `undef AXI_WPYLD_ID_RHS_M
`endif 

`ifdef AXI_WPYLD_ID_LHS_M
  `undef AXI_WPYLD_ID_LHS_M
`endif 

`ifdef AXI_WPYLD_ID_M
  `undef AXI_WPYLD_ID_M
`endif 

`ifdef AXI_WPYLD_ID_RHS_S
  `undef AXI_WPYLD_ID_RHS_S
`endif 

`ifdef AXI_WPYLD_ID_LHS_S
  `undef AXI_WPYLD_ID_LHS_S
`endif 

`ifdef AXI_WPYLD_ID_S
  `undef AXI_WPYLD_ID_S
`endif 

`ifdef AXI_BPYLD_RESP_RHS
  `undef AXI_BPYLD_RESP_RHS
`endif 

`ifdef AXI_BPYLD_RESP_LHS
  `undef AXI_BPYLD_RESP_LHS
`endif 

`ifdef AXI_BPYLD_RESP
  `undef AXI_BPYLD_RESP
`endif 

`ifdef AXI_BPYLD_ID_RHS_M
  `undef AXI_BPYLD_ID_RHS_M
`endif 

`ifdef AXI_BPYLD_ID_LHS_M
  `undef AXI_BPYLD_ID_LHS_M
`endif 

`ifdef AXI_BPYLD_ID_M
  `undef AXI_BPYLD_ID_M
`endif 

`ifdef AXI_BPYLD_ID_RHS_S
  `undef AXI_BPYLD_ID_RHS_S
`endif 

`ifdef AXI_BPYLD_ID_LHS_S
  `undef AXI_BPYLD_ID_LHS_S
`endif 

`ifdef AXI_BPYLD_ID_S
  `undef AXI_BPYLD_ID_S
`endif 

`ifdef AXI_QOSW
  `undef AXI_QOSW
`endif 

`ifdef IC_ADDR_SLICE_LHS
  `undef IC_ADDR_SLICE_LHS
`endif 

`ifdef MAX_APB_DATA_WIDTH
  `undef MAX_APB_DATA_WIDTH
`endif 

`ifdef REG_XCT_RATE_W
  `undef REG_XCT_RATE_W
`endif 

`ifdef REG_BURSTINESS_W
  `undef REG_BURSTINESS_W
`endif 

`ifdef REG_PEAK_RATE_W
  `undef REG_PEAK_RATE_W
`endif 

`ifdef APB_ADDR_WIDTH
  `undef APB_ADDR_WIDTH
`endif 

`ifdef AXI_ALSW
  `undef AXI_ALSW
`endif 

`ifdef AXI_ALDW
  `undef AXI_ALDW
`endif 

`ifdef AXI_ALBW
  `undef AXI_ALBW
`endif 

`ifdef AXI_REGIONW
  `undef AXI_REGIONW
`endif 

`ifdef PL_BUF_AW
  `undef PL_BUF_AW
`endif 

`ifdef PL_BUF_AR
  `undef PL_BUF_AR
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AW_M1
  `undef ACT_ID_BUF_POINTER_W_AW_M1
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AW_M1
  `undef LOG2_ACT_ID_BUF_POINTER_W_AW_M1
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AR_M1
  `undef ACT_ID_BUF_POINTER_W_AR_M1
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AR_M1
  `undef LOG2_ACT_ID_BUF_POINTER_W_AR_M1
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AW_M2
  `undef ACT_ID_BUF_POINTER_W_AW_M2
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AW_M2
  `undef LOG2_ACT_ID_BUF_POINTER_W_AW_M2
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AR_M2
  `undef ACT_ID_BUF_POINTER_W_AR_M2
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AR_M2
  `undef LOG2_ACT_ID_BUF_POINTER_W_AR_M2
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AW_M3
  `undef ACT_ID_BUF_POINTER_W_AW_M3
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AW_M3
  `undef LOG2_ACT_ID_BUF_POINTER_W_AW_M3
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AR_M3
  `undef ACT_ID_BUF_POINTER_W_AR_M3
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AR_M3
  `undef LOG2_ACT_ID_BUF_POINTER_W_AR_M3
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AW_M4
  `undef ACT_ID_BUF_POINTER_W_AW_M4
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AW_M4
  `undef LOG2_ACT_ID_BUF_POINTER_W_AW_M4
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AR_M4
  `undef ACT_ID_BUF_POINTER_W_AR_M4
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AR_M4
  `undef LOG2_ACT_ID_BUF_POINTER_W_AR_M4
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AW_M5
  `undef ACT_ID_BUF_POINTER_W_AW_M5
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AW_M5
  `undef LOG2_ACT_ID_BUF_POINTER_W_AW_M5
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AR_M5
  `undef ACT_ID_BUF_POINTER_W_AR_M5
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AR_M5
  `undef LOG2_ACT_ID_BUF_POINTER_W_AR_M5
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AW_M6
  `undef ACT_ID_BUF_POINTER_W_AW_M6
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AW_M6
  `undef LOG2_ACT_ID_BUF_POINTER_W_AW_M6
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AR_M6
  `undef ACT_ID_BUF_POINTER_W_AR_M6
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AR_M6
  `undef LOG2_ACT_ID_BUF_POINTER_W_AR_M6
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AW_M7
  `undef ACT_ID_BUF_POINTER_W_AW_M7
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AW_M7
  `undef LOG2_ACT_ID_BUF_POINTER_W_AW_M7
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AR_M7
  `undef ACT_ID_BUF_POINTER_W_AR_M7
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AR_M7
  `undef LOG2_ACT_ID_BUF_POINTER_W_AR_M7
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AW_M8
  `undef ACT_ID_BUF_POINTER_W_AW_M8
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AW_M8
  `undef LOG2_ACT_ID_BUF_POINTER_W_AW_M8
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AR_M8
  `undef ACT_ID_BUF_POINTER_W_AR_M8
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AR_M8
  `undef LOG2_ACT_ID_BUF_POINTER_W_AR_M8
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AW_M9
  `undef ACT_ID_BUF_POINTER_W_AW_M9
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AW_M9
  `undef LOG2_ACT_ID_BUF_POINTER_W_AW_M9
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AR_M9
  `undef ACT_ID_BUF_POINTER_W_AR_M9
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AR_M9
  `undef LOG2_ACT_ID_BUF_POINTER_W_AR_M9
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AW_M10
  `undef ACT_ID_BUF_POINTER_W_AW_M10
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AW_M10
  `undef LOG2_ACT_ID_BUF_POINTER_W_AW_M10
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AR_M10
  `undef ACT_ID_BUF_POINTER_W_AR_M10
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AR_M10
  `undef LOG2_ACT_ID_BUF_POINTER_W_AR_M10
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AW_M11
  `undef ACT_ID_BUF_POINTER_W_AW_M11
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AW_M11
  `undef LOG2_ACT_ID_BUF_POINTER_W_AW_M11
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AR_M11
  `undef ACT_ID_BUF_POINTER_W_AR_M11
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AR_M11
  `undef LOG2_ACT_ID_BUF_POINTER_W_AR_M11
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AW_M12
  `undef ACT_ID_BUF_POINTER_W_AW_M12
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AW_M12
  `undef LOG2_ACT_ID_BUF_POINTER_W_AW_M12
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AR_M12
  `undef ACT_ID_BUF_POINTER_W_AR_M12
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AR_M12
  `undef LOG2_ACT_ID_BUF_POINTER_W_AR_M12
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AW_M13
  `undef ACT_ID_BUF_POINTER_W_AW_M13
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AW_M13
  `undef LOG2_ACT_ID_BUF_POINTER_W_AW_M13
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AR_M13
  `undef ACT_ID_BUF_POINTER_W_AR_M13
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AR_M13
  `undef LOG2_ACT_ID_BUF_POINTER_W_AR_M13
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AW_M14
  `undef ACT_ID_BUF_POINTER_W_AW_M14
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AW_M14
  `undef LOG2_ACT_ID_BUF_POINTER_W_AW_M14
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AR_M14
  `undef ACT_ID_BUF_POINTER_W_AR_M14
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AR_M14
  `undef LOG2_ACT_ID_BUF_POINTER_W_AR_M14
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AW_M15
  `undef ACT_ID_BUF_POINTER_W_AW_M15
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AW_M15
  `undef LOG2_ACT_ID_BUF_POINTER_W_AW_M15
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AR_M15
  `undef ACT_ID_BUF_POINTER_W_AR_M15
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AR_M15
  `undef LOG2_ACT_ID_BUF_POINTER_W_AR_M15
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AW_M16
  `undef ACT_ID_BUF_POINTER_W_AW_M16
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AW_M16
  `undef LOG2_ACT_ID_BUF_POINTER_W_AW_M16
`endif 

`ifdef ACT_ID_BUF_POINTER_W_AR_M16
  `undef ACT_ID_BUF_POINTER_W_AR_M16
`endif 

`ifdef LOG2_ACT_ID_BUF_POINTER_W_AR_M16
  `undef LOG2_ACT_ID_BUF_POINTER_W_AR_M16
`endif 

`ifdef AXI_HAS_WID
  `undef AXI_HAS_WID
`endif 

`ifdef __GUARD__DW_AXI_BCM_PARAMS__VH__
  `undef __GUARD__DW_AXI_BCM_PARAMS__VH__
`endif 

`ifdef DW_AXI_RM_BCM00_AND
  `undef DW_AXI_RM_BCM00_AND
`endif 

`ifdef DW_AXI_RM_BCM00_ATPG_MX
  `undef DW_AXI_RM_BCM00_ATPG_MX
`endif 

`ifdef DW_AXI_RM_BCM00_CK_AND
  `undef DW_AXI_RM_BCM00_CK_AND
`endif 

`ifdef DW_AXI_RM_BCM00_CK_BUF
  `undef DW_AXI_RM_BCM00_CK_BUF
`endif 

`ifdef DW_AXI_RM_BCM00_CK_GT_LAT
  `undef DW_AXI_RM_BCM00_CK_GT_LAT
`endif 

`ifdef DW_AXI_RM_BCM00_CK_MX
  `undef DW_AXI_RM_BCM00_CK_MX
`endif 

`ifdef DW_AXI_RM_BCM00_CK_OR
  `undef DW_AXI_RM_BCM00_CK_OR
`endif 

`ifdef DW_AXI_RM_BCM00_MAJ
  `undef DW_AXI_RM_BCM00_MAJ
`endif 

`ifdef DW_AXI_RM_BCM00_MX
  `undef DW_AXI_RM_BCM00_MX
`endif 

`ifdef DW_AXI_RM_BCM00_OR
  `undef DW_AXI_RM_BCM00_OR
`endif 

`ifdef DW_AXI_RM_BCM01
  `undef DW_AXI_RM_BCM01
`endif 

`ifdef DW_AXI_RM_BCM02
  `undef DW_AXI_RM_BCM02
`endif 

`ifdef DW_AXI_RM_BCM03
  `undef DW_AXI_RM_BCM03
`endif 

`ifdef DW_AXI_RM_BCM04
  `undef DW_AXI_RM_BCM04
`endif 

`ifdef DW_AXI_RM_BCM05
  `undef DW_AXI_RM_BCM05
`endif 

`ifdef DW_AXI_RM_BCM05_ATV
  `undef DW_AXI_RM_BCM05_ATV
`endif 

`ifdef DW_AXI_RM_BCM05_CF
  `undef DW_AXI_RM_BCM05_CF
`endif 

`ifdef DW_AXI_RM_BCM05_EF
  `undef DW_AXI_RM_BCM05_EF
`endif 

`ifdef DW_AXI_RM_BCM05_EF_ATV
  `undef DW_AXI_RM_BCM05_EF_ATV
`endif 

`ifdef DW_AXI_RM_BCM06
  `undef DW_AXI_RM_BCM06
`endif 

`ifdef DW_AXI_RM_BCM06_ATV
  `undef DW_AXI_RM_BCM06_ATV
`endif 

`ifdef DW_AXI_RM_BCM07
  `undef DW_AXI_RM_BCM07
`endif 

`ifdef DW_AXI_RM_BCM07_ATV
  `undef DW_AXI_RM_BCM07_ATV
`endif 

`ifdef DW_AXI_RM_BCM07_EF
  `undef DW_AXI_RM_BCM07_EF
`endif 

`ifdef DW_AXI_RM_BCM07_EF_ATV
  `undef DW_AXI_RM_BCM07_EF_ATV
`endif 

`ifdef DW_AXI_RM_BCM07_EFES
  `undef DW_AXI_RM_BCM07_EFES
`endif 

`ifdef DW_AXI_RM_BCM07_RS
  `undef DW_AXI_RM_BCM07_RS
`endif 

`ifdef DW_AXI_RM_BCM08
  `undef DW_AXI_RM_BCM08
`endif 

`ifdef DW_AXI_RM_BCM09
  `undef DW_AXI_RM_BCM09
`endif 

`ifdef DW_AXI_RM_BCM09_DP
  `undef DW_AXI_RM_BCM09_DP
`endif 

`ifdef DW_AXI_RM_BCM09_ECC
  `undef DW_AXI_RM_BCM09_ECC
`endif 

`ifdef DW_AXI_RM_BCM10
  `undef DW_AXI_RM_BCM10
`endif 

`ifdef DW_AXI_RM_BCM11
  `undef DW_AXI_RM_BCM11
`endif 

`ifdef DW_AXI_RM_BCM12
  `undef DW_AXI_RM_BCM12
`endif 

`ifdef DW_AXI_RM_BCM14
  `undef DW_AXI_RM_BCM14
`endif 

`ifdef DW_AXI_RM_BCM15
  `undef DW_AXI_RM_BCM15
`endif 

`ifdef DW_AXI_RM_BCM16
  `undef DW_AXI_RM_BCM16
`endif 

`ifdef DW_AXI_RM_BCM17
  `undef DW_AXI_RM_BCM17
`endif 

`ifdef DW_AXI_RM_BCM18_GEN
  `undef DW_AXI_RM_BCM18_GEN
`endif 

`ifdef DW_AXI_RM_BCM18_MON
  `undef DW_AXI_RM_BCM18_MON
`endif 

`ifdef DW_AXI_RM_BCM18_PGEN
  `undef DW_AXI_RM_BCM18_PGEN
`endif 

`ifdef DW_AXI_RM_BCM18_PGENA
  `undef DW_AXI_RM_BCM18_PGENA
`endif 

`ifdef DW_AXI_RM_BCM18_PMON
  `undef DW_AXI_RM_BCM18_PMON
`endif 

`ifdef DW_AXI_RM_BCM18_RS
  `undef DW_AXI_RM_BCM18_RS
`endif 

`ifdef DW_AXI_RM_BCM19_INTR
  `undef DW_AXI_RM_BCM19_INTR
`endif 

`ifdef DW_AXI_RM_BCM19_TRGT
  `undef DW_AXI_RM_BCM19_TRGT
`endif 

`ifdef DW_AXI_RM_BCM21
  `undef DW_AXI_RM_BCM21
`endif 

`ifdef DW_AXI_RM_BCM21_ATV
  `undef DW_AXI_RM_BCM21_ATV
`endif 

`ifdef DW_AXI_RM_BCM21_NEO
  `undef DW_AXI_RM_BCM21_NEO
`endif 

`ifdef DW_AXI_RM_BCM21_TGL
  `undef DW_AXI_RM_BCM21_TGL
`endif 

`ifdef DW_AXI_RM_BCM22
  `undef DW_AXI_RM_BCM22
`endif 

`ifdef DW_AXI_RM_BCM22_ATV
  `undef DW_AXI_RM_BCM22_ATV
`endif 

`ifdef DW_AXI_RM_BCM23
  `undef DW_AXI_RM_BCM23
`endif 

`ifdef DW_AXI_RM_BCM23_ATV
  `undef DW_AXI_RM_BCM23_ATV
`endif 

`ifdef DW_AXI_RM_BCM23_C
  `undef DW_AXI_RM_BCM23_C
`endif 

`ifdef DW_AXI_RM_BCM24
  `undef DW_AXI_RM_BCM24
`endif 

`ifdef DW_AXI_RM_BCM24_AP
  `undef DW_AXI_RM_BCM24_AP
`endif 

`ifdef DW_AXI_RM_BCM25
  `undef DW_AXI_RM_BCM25
`endif 

`ifdef DW_AXI_RM_BCM25_ATV
  `undef DW_AXI_RM_BCM25_ATV
`endif 

`ifdef DW_AXI_RM_BCM25_C
  `undef DW_AXI_RM_BCM25_C
`endif 

`ifdef DW_AXI_RM_BCM26
  `undef DW_AXI_RM_BCM26
`endif 

`ifdef DW_AXI_RM_BCM26_ATV
  `undef DW_AXI_RM_BCM26_ATV
`endif 

`ifdef DW_AXI_RM_BCM27
  `undef DW_AXI_RM_BCM27
`endif 

`ifdef DW_AXI_RM_BCM28
  `undef DW_AXI_RM_BCM28
`endif 

`ifdef DW_AXI_RM_BCM29
  `undef DW_AXI_RM_BCM29
`endif 

`ifdef DW_AXI_RM_BCM31_P2D_FIFOMEM
  `undef DW_AXI_RM_BCM31_P2D_FIFOMEM
`endif 

`ifdef DW_AXI_RM_BCM31_P2D_RD
  `undef DW_AXI_RM_BCM31_P2D_RD
`endif 

`ifdef DW_AXI_RM_BCM31_P2D_WR
  `undef DW_AXI_RM_BCM31_P2D_WR
`endif 

`ifdef DW_AXI_RM_BCM32_A
  `undef DW_AXI_RM_BCM32_A
`endif 

`ifdef DW_AXI_RM_BCM32_C
  `undef DW_AXI_RM_BCM32_C
`endif 

`ifdef DW_AXI_RM_BCM33_63_7_64_0
  `undef DW_AXI_RM_BCM33_63_7_64_0
`endif 

`ifdef DW_AXI_RM_BCM35
  `undef DW_AXI_RM_BCM35
`endif 

`ifdef DW_AXI_RM_BCM35_T
  `undef DW_AXI_RM_BCM35_T
`endif 

`ifdef DW_AXI_RM_BCM36
  `undef DW_AXI_RM_BCM36
`endif 

`ifdef DW_AXI_RM_BCM36_ACK
  `undef DW_AXI_RM_BCM36_ACK
`endif 

`ifdef DW_AXI_RM_BCM36_NHS
  `undef DW_AXI_RM_BCM36_NHS
`endif 

`ifdef DW_AXI_RM_BCM36_TGL
  `undef DW_AXI_RM_BCM36_TGL
`endif 

`ifdef DW_AXI_RM_BCM36_TGL_DO
  `undef DW_AXI_RM_BCM36_TGL_DO
`endif 

`ifdef DW_AXI_RM_BCM36_TGL_PLS
  `undef DW_AXI_RM_BCM36_TGL_PLS
`endif 

`ifdef DW_AXI_RM_BCM36_TGL_PLS_DO
  `undef DW_AXI_RM_BCM36_TGL_PLS_DO
`endif 

`ifdef DW_AXI_RM_BCM37
  `undef DW_AXI_RM_BCM37
`endif 

`ifdef DW_AXI_RM_BCM38
  `undef DW_AXI_RM_BCM38
`endif 

`ifdef DW_AXI_RM_BCM38_ADP
  `undef DW_AXI_RM_BCM38_ADP
`endif 

`ifdef DW_AXI_RM_BCM38_AP
  `undef DW_AXI_RM_BCM38_AP
`endif 

`ifdef DW_AXI_RM_BCM38_ECC
  `undef DW_AXI_RM_BCM38_ECC
`endif 

`ifdef DW_AXI_RM_BCM39
  `undef DW_AXI_RM_BCM39
`endif 

`ifdef DW_AXI_RM_BCM40
  `undef DW_AXI_RM_BCM40
`endif 

`ifdef DW_AXI_RM_BCM41
  `undef DW_AXI_RM_BCM41
`endif 

`ifdef DW_AXI_RM_BCM41_NEO
  `undef DW_AXI_RM_BCM41_NEO
`endif 

`ifdef DW_AXI_RM_BCM43
  `undef DW_AXI_RM_BCM43
`endif 

`ifdef DW_AXI_RM_BCM43_NRO
  `undef DW_AXI_RM_BCM43_NRO
`endif 

`ifdef DW_AXI_RM_BCM44
  `undef DW_AXI_RM_BCM44
`endif 

`ifdef DW_AXI_RM_BCM44_NRO
  `undef DW_AXI_RM_BCM44_NRO
`endif 

`ifdef DW_AXI_RM_BCM45_GN_D_A
  `undef DW_AXI_RM_BCM45_GN_D_A
`endif 

`ifdef DW_AXI_RM_BCM45_GN_D_AA
  `undef DW_AXI_RM_BCM45_GN_D_AA
`endif 

`ifdef DW_AXI_RM_BCM45_GN_D_B
  `undef DW_AXI_RM_BCM45_GN_D_B
`endif 

`ifdef DW_AXI_RM_BCM45_GN_D_C
  `undef DW_AXI_RM_BCM45_GN_D_C
`endif 

`ifdef DW_AXI_RM_BCM45_GN_D_D
  `undef DW_AXI_RM_BCM45_GN_D_D
`endif 

`ifdef DW_AXI_RM_BCM45_GN_D_E
  `undef DW_AXI_RM_BCM45_GN_D_E
`endif 

`ifdef DW_AXI_RM_BCM45_GN_D_F
  `undef DW_AXI_RM_BCM45_GN_D_F
`endif 

`ifdef DW_AXI_RM_BCM45_MN_D_A
  `undef DW_AXI_RM_BCM45_MN_D_A
`endif 

`ifdef DW_AXI_RM_BCM45_MN_D_AA
  `undef DW_AXI_RM_BCM45_MN_D_AA
`endif 

`ifdef DW_AXI_RM_BCM45_MN_D_B
  `undef DW_AXI_RM_BCM45_MN_D_B
`endif 

`ifdef DW_AXI_RM_BCM45_MN_D_C
  `undef DW_AXI_RM_BCM45_MN_D_C
`endif 

`ifdef DW_AXI_RM_BCM45_MN_D_D
  `undef DW_AXI_RM_BCM45_MN_D_D
`endif 

`ifdef DW_AXI_RM_BCM45_MN_D_E
  `undef DW_AXI_RM_BCM45_MN_D_E
`endif 

`ifdef DW_AXI_RM_BCM45_MN_D_F
  `undef DW_AXI_RM_BCM45_MN_D_F
`endif 

`ifdef DW_AXI_RM_BCM46_A
  `undef DW_AXI_RM_BCM46_A
`endif 

`ifdef DW_AXI_RM_BCM46_AA
  `undef DW_AXI_RM_BCM46_AA
`endif 

`ifdef DW_AXI_RM_BCM46_B
  `undef DW_AXI_RM_BCM46_B
`endif 

`ifdef DW_AXI_RM_BCM46_B_32A
  `undef DW_AXI_RM_BCM46_B_32A
`endif 

`ifdef DW_AXI_RM_BCM46_C
  `undef DW_AXI_RM_BCM46_C
`endif 

`ifdef DW_AXI_RM_BCM46_C_64A
  `undef DW_AXI_RM_BCM46_C_64A
`endif 

`ifdef DW_AXI_RM_BCM46_D
  `undef DW_AXI_RM_BCM46_D
`endif 

`ifdef DW_AXI_RM_BCM46_D_128A
  `undef DW_AXI_RM_BCM46_D_128A
`endif 

`ifdef DW_AXI_RM_BCM46_E
  `undef DW_AXI_RM_BCM46_E
`endif 

`ifdef DW_AXI_RM_BCM46_F
  `undef DW_AXI_RM_BCM46_F
`endif 

`ifdef DW_AXI_RM_BCM46_X
  `undef DW_AXI_RM_BCM46_X
`endif 

`ifdef DW_AXI_RM_BCM47
  `undef DW_AXI_RM_BCM47
`endif 

`ifdef DW_AXI_RM_BCM48
  `undef DW_AXI_RM_BCM48
`endif 

`ifdef DW_AXI_RM_BCM48_DM
  `undef DW_AXI_RM_BCM48_DM
`endif 

`ifdef DW_AXI_RM_BCM48_SV
  `undef DW_AXI_RM_BCM48_SV
`endif 

`ifdef DW_AXI_RM_BCM49
  `undef DW_AXI_RM_BCM49
`endif 

`ifdef DW_AXI_RM_BCM49_SV
  `undef DW_AXI_RM_BCM49_SV
`endif 

`ifdef DW_AXI_RM_BCM50
  `undef DW_AXI_RM_BCM50
`endif 

`ifdef DW_AXI_RM_BCM51
  `undef DW_AXI_RM_BCM51
`endif 

`ifdef DW_AXI_RM_BCM52
  `undef DW_AXI_RM_BCM52
`endif 

`ifdef DW_AXI_RM_BCM53
  `undef DW_AXI_RM_BCM53
`endif 

`ifdef DW_AXI_RM_BCM54
  `undef DW_AXI_RM_BCM54
`endif 

`ifdef DW_AXI_RM_BCM55
  `undef DW_AXI_RM_BCM55
`endif 

`ifdef DW_AXI_RM_BCM55_C
  `undef DW_AXI_RM_BCM55_C
`endif 

`ifdef DW_AXI_RM_BCM56
  `undef DW_AXI_RM_BCM56
`endif 

`ifdef DW_AXI_RM_BCM57
  `undef DW_AXI_RM_BCM57
`endif 

`ifdef DW_AXI_RM_BCM57_ATV
  `undef DW_AXI_RM_BCM57_ATV
`endif 

`ifdef DW_AXI_RM_BCM58
  `undef DW_AXI_RM_BCM58
`endif 

`ifdef DW_AXI_RM_BCM58_ATV
  `undef DW_AXI_RM_BCM58_ATV
`endif 

`ifdef DW_AXI_RM_BCM59
  `undef DW_AXI_RM_BCM59
`endif 

`ifdef DW_AXI_RM_BCM60
  `undef DW_AXI_RM_BCM60
`endif 

`ifdef DW_AXI_RM_BCM62
  `undef DW_AXI_RM_BCM62
`endif 

`ifdef DW_AXI_RM_BCM63
  `undef DW_AXI_RM_BCM63
`endif 

`ifdef DW_AXI_RM_BCM64
  `undef DW_AXI_RM_BCM64
`endif 

`ifdef DW_AXI_RM_BCM64_TD
  `undef DW_AXI_RM_BCM64_TD
`endif 

`ifdef DW_AXI_RM_BCM65
  `undef DW_AXI_RM_BCM65
`endif 

`ifdef DW_AXI_RM_BCM65_ATV
  `undef DW_AXI_RM_BCM65_ATV
`endif 

`ifdef DW_AXI_RM_BCM65_TD
  `undef DW_AXI_RM_BCM65_TD
`endif 

`ifdef DW_AXI_RM_BCM66
  `undef DW_AXI_RM_BCM66
`endif 

`ifdef DW_AXI_RM_BCM66_ATV
  `undef DW_AXI_RM_BCM66_ATV
`endif 

`ifdef DW_AXI_RM_BCM66_DMS
  `undef DW_AXI_RM_BCM66_DMS
`endif 

`ifdef DW_AXI_RM_BCM66_DMS_ATV
  `undef DW_AXI_RM_BCM66_DMS_ATV
`endif 

`ifdef DW_AXI_RM_BCM66_EFES
  `undef DW_AXI_RM_BCM66_EFES
`endif 

`ifdef DW_AXI_RM_BCM66_PR
  `undef DW_AXI_RM_BCM66_PR
`endif 

`ifdef DW_AXI_RM_BCM66_WAE
  `undef DW_AXI_RM_BCM66_WAE
`endif 

`ifdef DW_AXI_RM_BCM66_WAE_ATV
  `undef DW_AXI_RM_BCM66_WAE_ATV
`endif 

`ifdef DW_AXI_RM_BCM68_63_7_0
  `undef DW_AXI_RM_BCM68_63_7_0
`endif 

`ifdef DW_AXI_RM_BCM69_63_7_0
  `undef DW_AXI_RM_BCM69_63_7_0
`endif 

`ifdef DW_AXI_RM_BCM70_63_7_0_0
  `undef DW_AXI_RM_BCM70_63_7_0_0
`endif 

`ifdef DW_AXI_RM_BCM71
  `undef DW_AXI_RM_BCM71
`endif 

`ifdef DW_AXI_RM_BCM72
  `undef DW_AXI_RM_BCM72
`endif 

`ifdef DW_AXI_RM_BCM74
  `undef DW_AXI_RM_BCM74
`endif 

`ifdef DW_AXI_RM_BCM76
  `undef DW_AXI_RM_BCM76
`endif 

`ifdef DW_AXI_RM_BCM77
  `undef DW_AXI_RM_BCM77
`endif 

`ifdef DW_AXI_RM_BCM78
  `undef DW_AXI_RM_BCM78
`endif 

`ifdef DW_AXI_RM_BCM79
  `undef DW_AXI_RM_BCM79
`endif 

`ifdef DW_AXI_RM_BCM79_MO
  `undef DW_AXI_RM_BCM79_MO
`endif 

`ifdef DW_AXI_RM_BCM83_GEN
  `undef DW_AXI_RM_BCM83_GEN
`endif 

`ifdef DW_AXI_RM_BCM84_MON
  `undef DW_AXI_RM_BCM84_MON
`endif 

`ifdef DW_AXI_RM_BCM85
  `undef DW_AXI_RM_BCM85
`endif 

`ifdef DW_AXI_RM_BCM86
  `undef DW_AXI_RM_BCM86
`endif 

`ifdef DW_AXI_RM_BCM87
  `undef DW_AXI_RM_BCM87
`endif 

`ifdef DW_AXI_RM_BCM90
  `undef DW_AXI_RM_BCM90
`endif 

`ifdef DW_AXI_RM_BCM91
  `undef DW_AXI_RM_BCM91
`endif 

`ifdef DW_AXI_RM_BCM92
  `undef DW_AXI_RM_BCM92
`endif 

`ifdef DW_AXI_RM_BCM92_AD
  `undef DW_AXI_RM_BCM92_AD
`endif 

`ifdef DW_AXI_RM_BCM92_AD_DO
  `undef DW_AXI_RM_BCM92_AD_DO
`endif 

`ifdef DW_AXI_RM_BCM92_RD
  `undef DW_AXI_RM_BCM92_RD
`endif 

`ifdef DW_AXI_RM_BCM92_RD_AD
  `undef DW_AXI_RM_BCM92_RD_AD
`endif 

`ifdef DW_AXI_RM_BCM92_RD_AD_DO
  `undef DW_AXI_RM_BCM92_RD_AD_DO
`endif 

`ifdef DW_AXI_RM_BCM92_RD_DO
  `undef DW_AXI_RM_BCM92_RD_DO
`endif 

`ifdef DW_AXI_RM_BCM93
  `undef DW_AXI_RM_BCM93
`endif 

`ifdef DW_AXI_RM_BCM93_NDSVA
  `undef DW_AXI_RM_BCM93_NDSVA
`endif 

`ifdef DW_AXI_RM_BCM94
  `undef DW_AXI_RM_BCM94
`endif 

`ifdef DW_AXI_RM_BCM95
  `undef DW_AXI_RM_BCM95
`endif 

`ifdef DW_AXI_RM_BCM95_E
  `undef DW_AXI_RM_BCM95_E
`endif 

`ifdef DW_AXI_RM_BCM95_I
  `undef DW_AXI_RM_BCM95_I
`endif 

`ifdef DW_AXI_RM_BCM95_IE
  `undef DW_AXI_RM_BCM95_IE
`endif 

`ifdef DW_AXI_RM_BCM95_NE
  `undef DW_AXI_RM_BCM95_NE
`endif 

`ifdef DW_AXI_RM_BCM95_NE_E
  `undef DW_AXI_RM_BCM95_NE_E
`endif 

`ifdef DW_AXI_RM_BCM95_NE_I
  `undef DW_AXI_RM_BCM95_NE_I
`endif 

`ifdef DW_AXI_RM_BCM95_NE_IE
  `undef DW_AXI_RM_BCM95_NE_IE
`endif 

`ifdef DW_AXI_RM_BCM98
  `undef DW_AXI_RM_BCM98
`endif 

`ifdef DW_AXI_RM_BCM99
  `undef DW_AXI_RM_BCM99
`endif 

`ifdef DW_AXI_RM_BCM99_3
  `undef DW_AXI_RM_BCM99_3
`endif 

`ifdef DW_AXI_RM_BCM99_4
  `undef DW_AXI_RM_BCM99_4
`endif 

`ifdef DW_AXI_RM_BCM99_N
  `undef DW_AXI_RM_BCM99_N
`endif 

`ifdef DW_AXI_RM_BVM01
  `undef DW_AXI_RM_BVM01
`endif 

`ifdef DW_AXI_RM_BVM02
  `undef DW_AXI_RM_BVM02
`endif 

`ifdef DW_AXI_RM_SVA01
  `undef DW_AXI_RM_SVA01
`endif 

`ifdef DW_AXI_RM_SVA02
  `undef DW_AXI_RM_SVA02
`endif 

`ifdef DW_AXI_RM_SVA03
  `undef DW_AXI_RM_SVA03
`endif 

`ifdef DW_AXI_RM_SVA04
  `undef DW_AXI_RM_SVA04
`endif 

`ifdef DW_AXI_RM_SVA05
  `undef DW_AXI_RM_SVA05
`endif 

`ifdef DW_AXI_RM_SVA06
  `undef DW_AXI_RM_SVA06
`endif 

`ifdef DW_AXI_RM_SVA07
  `undef DW_AXI_RM_SVA07
`endif 

`ifdef DW_AXI_RM_SVA08
  `undef DW_AXI_RM_SVA08
`endif 

`ifdef DW_AXI_RM_SVA09
  `undef DW_AXI_RM_SVA09
`endif 

`ifdef DW_AXI_RM_SVA10
  `undef DW_AXI_RM_SVA10
`endif 

`ifdef DW_AXI_RM_SVA11
  `undef DW_AXI_RM_SVA11
`endif 

`ifdef DW_AXI_RM_SVA12_A
  `undef DW_AXI_RM_SVA12_A
`endif 

`ifdef DW_AXI_RM_SVA12_B
  `undef DW_AXI_RM_SVA12_B
`endif 

`ifdef DW_AXI_RM_SVA12_C
  `undef DW_AXI_RM_SVA12_C
`endif 

`ifdef DW_AXI_RM_SVA99
  `undef DW_AXI_RM_SVA99
`endif 

`ifdef __GUARD__DW_AXI_ALL_INCLUDES__VH__
  `undef __GUARD__DW_AXI_ALL_INCLUDES__VH__
`endif 

`ifdef DW_HOLD_MUX_DELAY
  `undef DW_HOLD_MUX_DELAY
`endif 

`ifdef DW_SETUP_MUX_DELAY
  `undef DW_SETUP_MUX_DELAY
`endif 

`ifdef cb_dummy_parameter_definition
  `undef cb_dummy_parameter_definition
`endif 

